magic
tech sky130A
magscale 1 2
timestamp 1739996415
<< error_s >>
rect 9030 -840 10068 -554
rect 9030 -1374 9316 -840
rect 9520 -990 9578 -984
rect 9520 -1024 9532 -990
rect 9520 -1030 9578 -1024
rect 9527 -1152 9571 -1062
rect 9520 -1190 9578 -1184
rect 9520 -1224 9532 -1190
rect 9520 -1230 9578 -1224
rect 9782 -1374 10068 -840
rect 9030 -1660 10068 -1374
use sky130_fd_bs_flash__special_sonosfet_star_EA7MKQ  X1
timestamp 1739996415
transform 1 0 9549 0 1 -1107
box -519 -553 519 553
use charge_pump_neg_nmos  x2 ../charge_pump_neg_nmos
timestamp 1739484054
transform 1 0 10614 0 1 18680
box -4288 -1488 12990 4458
use charge_pump  x3 ../charge_pump
timestamp 1739252499
transform 1 0 10730 0 1 11954
box -4288 -1488 12990 4458
use vprog_controller  x4 ../vprog_controller
timestamp 1738900598
transform 1 0 23018 0 1 22946
box 1324 -4282 4846 -1260
use inverter  x5 ../inverter
timestamp 1739087840
transform 1 0 36328 0 1 16172
box 0 -620 992 638
use inverter  x6
timestamp 1739087840
transform 1 0 30140 0 1 14922
box 0 -620 992 638
use vprog_controller  x7
timestamp 1738900598
transform 1 0 22738 0 1 17336
box 1324 -4282 4846 -1260
use sky130_fd_pr__pfet_g5v0d10v5_VPAE37  XM1
timestamp 1739996415
transform 1 0 15058 0 1 2187
box -2258 -347 2258 347
use sky130_fd_pr__pfet_g5v0d10v5_VPAE37  XM2
timestamp 1739996415
transform 1 0 15058 0 1 1493
box -2258 -347 2258 347
use sky130_fd_pr__pfet_g5v0d10v5_GJ3XY6  XM3
timestamp 1739996415
transform 1 0 14058 0 1 799
box -1258 -347 1258 347
use sky130_fd_pr__pfet_g5v0d10v5_VPAE37  XM4
timestamp 1739996415
transform 1 0 33614 0 1 16325
box -2258 -347 2258 347
use sky130_fd_pr__nfet_g5v0d10v5_9UU773  XM5
timestamp 1739996415
transform 1 0 8472 0 1 970
box -278 -758 278 758
use sky130_fd_pr__nfet_g5v0d10v5_HQS8YU  XM8
timestamp 1739996415
transform 1 0 10566 0 1 528
box -278 -458 278 458
<< end >>
