** sch_path: /home/amedcalf/projects/tt10-sonos-flash-party/xschem/vprog_controller_tb.sch
**.subckt vprog_controller_tb
V1 VPRGNEG GND -3.7
V3 VDPWR GND 1.8
x1 pos_en neg_en vout VDPWR net1 VPRGPOS VPRGNEG vprog_controller
V4 neg_en GND PULSE(0 1.8 4u 0 0 1u 1s)
V5 pos_en GND PULSE(0 1.8 2u 0 0 1u 1s)
V2 VPRGPOS GND 6.7
V6 net1 GND 0
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/amedcalf/open-asic/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt
.include ../../spice/vprog_controller/pex/vprog_controller.spice




.option savecurrents
.tran 1n 10u
.save all

.control
run
remzerovec
write vprog_controller_tb.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
