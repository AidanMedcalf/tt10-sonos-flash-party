* NGSPICE file created from tt_um_sonos_flash_party.ext - technology: sky130A

.subckt tt_um_sonos_flash_party clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VDPWR VGND VAPWR
X0 flash_0.x7.VPRGNEG VGND.t51 sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X1 flash_0.x7.VPRGPOS.t25 flash_0.x7.pos_mid_b.t3 flash_0.x7.vintp flash_0.x7.VPRGPOS.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X2 flash_0.x2.clkb.t0 flash_0.x2.clkinb VAPWR.t12 VAPWR.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X3 flash_0.x7.VPRGPOS.t26 flash_0.x7.pos_mid flash_0.x7.pos_mid_b.t1 flash_0.x7.VPRGPOS.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X4 flash_0.x3.clkinb clk.t0 VAPWR.t1 VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X5 flash_0.x7.VPRGPOS.t7 flash_0.x4.pos_mid flash_0.x4.pos_mid_b.t1 flash_0.x7.VPRGPOS.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X6 VGND.t9 ui_in[1].t0 flash_0.x4.neg_en_b.t2 VGND.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X7 flash_0.x4.dcgint.t11 flash_0.x4.neg_mid_b.t7 flash_0.x4.VOUT.t8 flash_0.x4.dcgint.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X8 flash_0.x7.pos_mid_b.t2 ui_in[1].t1 VGND.t61 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X9 flash_0.x7.pos_mid flash_0.x7.pos_en_b.t4 VGND.t24 VGND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X10 VDPWR.t40 ui_in[1].t2 flash_0.x4.neg_mid VDPWR.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X11 ua[0].t3 VGND.t49 VGND.t50 ua[0].t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=10
X12 VDPWR.t56 flash_0.x7.neg_en_b.t4 flash_0.x7.neg_mid_b.t5 VDPWR.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X13 VDPWR.t52 flash_0.x7.neg_en_b.t5 flash_0.x7.neg_mid_b.t4 VDPWR.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X14 flash_0.x5.A.t3 flash_0.x6.Y VDPWR.t54 VDPWR.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
X15 flash_0.x7.vintp flash_0.x7.pos_mid_b.t4 flash_0.x7.VPRGPOS.t23 flash_0.x7.VPRGPOS.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X16 flash_0.x7.neg_mid ui_in[0].t0 VDPWR.t18 VDPWR.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X17 flash_0.x4.neg_mid_b.t0 flash_0.x4.neg_mid flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=1
X18 flash_0.x2.clkina flash_0.x2.clkinb VAPWR.t10 VAPWR.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X19 flash_0.x4.neg_mid_b.t5 flash_0.x4.neg_en_b.t4 VDPWR.t51 VDPWR.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X20 flash_0.x7.pos_mid_b.t0 ui_in[1].t3 VGND.t35 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X21 flash_0.x7.pos_mid flash_0.x7.pos_en_b.t4 VGND.t23 VGND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X22 flash_0.x4.dcgint.t10 flash_0.x4.neg_mid_b.t8 flash_0.x4.VOUT.t10 flash_0.x4.dcgint.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X23 a_9352_28387# flash_0.x4.VOUT.t14 a_7463_28281# flash_0.x7.VOUT.t0 sky130_fd_bs_flash__special_sonosfet_star ad=0.13725 pd=1.51 as=0.13725 ps=1.51 w=0.45 l=0.22
X24 VGND.t18 ui_in[1].t4 flash_0.x7.pos_mid_b VGND.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X25 VGND.t5 ui_in[0].t1 flash_0.x4.pos_mid_b VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X26 flash_0.x7.VPRGNEG flash_0.x4.neg_mid_b.t9 flash_0.x4.neg_mid flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.145 ps=1.58 w=0.5 l=1
X27 flash_0.x4.vintp VDPWR.t58 flash_0.x4.VOUT.t2 flash_0.x7.VPRGPOS.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X28 VDPWR.t38 ui_in[1].t5 flash_0.x4.neg_en_b.t3 VDPWR.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X29 flash_0.x4.VOUT.t0 VDPWR.t59 a_16296_28578# flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X30 VDPWR.t41 flash_0.x7.neg_en_b.t6 flash_0.x7.neg_mid_b.t3 VDPWR.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X31 w_7728_24730.t1 ua[0].t0 ua[0].t1 w_7728_24730.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
X32 flash_0.x3.stage1 VAPWR.t2 VAPWR.t4 VAPWR.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X33 flash_0.x4.VOUT.t5 VDPWR.t60 flash_0.x4.vintp flash_0.x7.VPRGPOS.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X34 flash_0.x7.neg_en_b.t1 ui_in[0].t2 VGND.t1 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X35 flash_0.x7.pos_en_b.t3 ui_in[1].t6 VGND.t47 VGND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X36 VGND.t60 ui_in[1].t7 flash_0.x7.pos_mid_b VGND.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X37 flash_0.x3.clka.t0 flash_0.x3.clkina VAPWR.t8 VAPWR.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X38 VGND.t68 ui_in[0].t3 flash_0.x4.pos_mid_b VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X39 flash_0.x3.clkb.t1 flash_0.x3.clkinb VGND.t59 VGND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X40 flash_0.x4.vintp flash_0.x4.pos_mid_b.t3 flash_0.x7.VPRGPOS.t10 flash_0.x7.VPRGPOS.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X41 flash_0.x4.VOUT.t4 VDPWR.t61 a_16296_28578# flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X42 flash_0.x4.dcgint.t2 flash_0.x4.pos_en_b.t4 VGND.t33 VGND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X43 flash_0.x7.VPRGPOS.t4 flash_0.x4.pos_mid_b.t4 flash_0.x4.vintp flash_0.x7.VPRGPOS.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X44 flash_0.x6.Y.t0 ui_in[2].t0 VGND.t15 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X45 flash_0.x7.VOUT.t8 VDPWR.t62 flash_0.x7.vintp flash_0.x7.VPRGPOS.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X46 flash_0.x2.clka.t1 flash_0.x2.clkina VGND.t63 VGND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X47 flash_0.x3.clkb flash_0.x3.stage2 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X48 VGND.t34 ui_in[1].t8 flash_0.x7.pos_en_b.t2 VGND.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X49 VGND.t48 ui_in[0].t4 flash_0.x4.pos_en_b.t3 VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X50 VDPWR.t50 flash_0.x4.neg_en_b.t5 flash_0.x4.neg_mid_b.t1 VDPWR.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X51 flash_0.x7.neg_en_b.t2 ui_in[0].t5 VDPWR.t20 VDPWR.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=3
X52 flash_0.x7.pos_en_b.t1 ui_in[1].t9 VDPWR.t36 VDPWR.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X53 flash_0.x4.dcgint.t1 flash_0.x4.pos_en_b.t4 VGND.t31 VGND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X54 VDPWR.t34 ui_in[1].t10 flash_0.x4.neg_mid VDPWR.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X55 a_16296_28578# flash_0.x4.neg_mid_b.t10 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X56 flash_0.x4.neg_mid_b.t4 flash_0.x4.neg_en_b.t6 VDPWR.t49 VDPWR.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X57 flash_0.x7.VPRGPOS.t22 flash_0.x7.pos_mid_b.t5 flash_0.x7.vintp flash_0.x7.VPRGPOS.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X58 flash_0.x7.neg_mid ui_in[0].t6 VDPWR.t9 VDPWR.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X59 flash_0.x4.neg_mid_b.t6 flash_0.x4.neg_en_b.t7 VDPWR.t48 VDPWR.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X60 flash_0.x4.dcgint.t8 flash_0.x4.neg_mid_b.t11 flash_0.x4.VOUT.t11 flash_0.x4.dcgint.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X61 flash_0.x7.VPRGPOS.t29 w_7728_24730.t2 w_7728_24730.t3 flash_0.x7.VPRGPOS.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
X62 VDPWR.t32 ui_in[1].t11 flash_0.x7.pos_en_b.t0 VDPWR.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X63 flash_0.x3.clkinb clk.t1 VGND.t11 VGND.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X64 VDPWR.t7 ui_in[0].t7 flash_0.x4.pos_en_b.t1 VDPWR.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X65 flash_0.x2.clkina flash_0.x2.clkinb VGND.t55 VGND.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X66 flash_0.x3.clka flash_0.x3.stage1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X67 a_16296_28578# flash_0.x4.neg_mid_b.t10 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X68 flash_0.x4.dcgint.t0 flash_0.x4.pos_en_b.t4 VGND.t29 VGND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X69 flash_0.x4.VOUT.t9 flash_0.x4.neg_mid_b.t12 flash_0.x4.dcgint.t7 flash_0.x4.dcgint.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X70 flash_0.x4.dcgint.t6 flash_0.x4.neg_mid_b.t13 flash_0.x4.VOUT.t7 flash_0.x4.dcgint.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X71 flash_0.x4.vintp VDPWR.t63 flash_0.x4.VOUT.t1 flash_0.x7.VPRGPOS.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X72 a_7463_28281# ui_in[2].t1 VGND.t67 VGND.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X73 flash_0.x7.neg_mid ui_in[0].t8 VDPWR.t57 VDPWR.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X74 flash_0.x7.dcgint.t8 flash_0.x7.neg_mid_b.t7 flash_0.x7.VOUT.t14 flash_0.x7.dcgint.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X75 VDPWR.t43 ui_in[0].t9 flash_0.x7.neg_mid VDPWR.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X76 uo_out[0].t0 flash_0.x5.A.t4 VDPWR.t45 VDPWR.t44 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X77 VDPWR.t3 ui_in[0].t10 flash_0.x7.neg_mid VDPWR.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X78 flash_0.x4.VOUT.t12 VDPWR.t64 flash_0.x4.vintp flash_0.x7.VPRGPOS.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X79 flash_0.x3.stage2 flash_0.x3.stage1 flash_0.x3.stage1 flash_0.x3.stage1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X80 flash_0.x2.clkinb clk.t2 VAPWR.t6 VAPWR.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X81 flash_0.x4.VOUT.t6 flash_0.x4.neg_mid_b.t14 flash_0.x4.dcgint.t4 flash_0.x4.dcgint.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X82 flash_0.x7.neg_mid_b.t6 flash_0.x7.neg_mid flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=1
X83 flash_0.x4.vintp flash_0.x4.pos_mid_b.t5 flash_0.x7.VPRGPOS.t5 flash_0.x7.VPRGPOS.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X84 VGND.t38 flash_0.x7.pos_en_b.t5 flash_0.x7.pos_mid VGND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X85 flash_0.x7.dcgint.t7 flash_0.x7.neg_mid_b.t8 flash_0.x7.VOUT.t9 flash_0.x7.dcgint.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X86 flash_0.x3.clkb.t0 flash_0.x3.clkinb VAPWR.t15 VAPWR.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X87 flash_0.x7.vintp VDPWR.t65 flash_0.x7.VOUT.t7 flash_0.x7.VPRGPOS.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X88 flash_0.x7.VOUT.t2 VDPWR.t66 a_20416_28577# flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X89 flash_0.x4.vintp VDPWR.t67 flash_0.x4.VOUT.t13 flash_0.x7.VPRGPOS.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X90 flash_0.x7.VPRGPOS.t32 flash_0.x4.pos_mid_b.t6 flash_0.x4.vintp flash_0.x7.VPRGPOS.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X91 flash_0.x2.clkb flash_0.x2.stage2 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X92 flash_0.x2.stage1 flash_0.x2.stage1 VGND.t19 flash_0.x2.stage1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X93 flash_0.x7.VPRGPOS.t11 flash_0.x3.stage2 flash_0.x3.stage2 flash_0.x3.stage2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X94 VGND.t37 flash_0.x7.pos_en_b.t5 flash_0.x7.pos_mid VGND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X95 flash_0.x4.pos_mid_b.t0 ui_in[0].t11 VGND.t13 VGND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X96 flash_0.x4.pos_mid flash_0.x4.pos_en_b.t5 VGND.t65 VGND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X97 flash_0.x2.clkb.t1 flash_0.x2.clkinb VGND.t53 VGND.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X98 flash_0.x3.clkina flash_0.x3.clkinb VAPWR.t14 VAPWR.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X99 flash_0.x7.vintp flash_0.x7.pos_mid_b.t6 flash_0.x7.VPRGPOS.t21 flash_0.x7.VPRGPOS.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X100 VDPWR.t47 flash_0.x4.neg_en_b.t8 flash_0.x4.neg_mid_b.t2 VDPWR.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X101 flash_0.x7.VOUT.t1 VDPWR.t68 a_20416_28577# flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X102 flash_0.x4.vintp flash_0.x4.pos_mid_b.t7 flash_0.x7.VPRGPOS.t16 flash_0.x7.VPRGPOS.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X103 flash_0.x7.dcgint.t11 flash_0.x7.pos_en_b.t6 VGND.t44 VGND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X104 a_20416_28577# flash_0.x7.neg_mid_b.t9 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X105 flash_0.x2.clka.t0 flash_0.x2.clkina VAPWR.t16 VAPWR.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X106 VGND.t70 ui_in[0].t12 flash_0.x7.neg_en_b.t3 VGND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X107 flash_0.x7.neg_mid_b.t2 flash_0.x7.neg_en_b.t7 VDPWR.t5 VDPWR.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X108 flash_0.x4.pos_mid_b.t2 ui_in[0].t13 VGND.t27 VGND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X109 flash_0.x4.neg_mid ui_in[1].t12 VDPWR.t30 VDPWR.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X110 flash_0.x4.pos_mid flash_0.x4.pos_en_b.t5 VGND.t64 VGND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X111 VDPWR.t28 ui_in[1].t13 flash_0.x4.neg_mid VDPWR.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X112 flash_0.x2.clka flash_0.x2.stage1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X113 flash_0.x7.VPRGPOS VGND.t69 sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X114 VDPWR.t46 flash_0.x4.neg_en_b.t9 flash_0.x4.neg_mid_b.t3 VDPWR.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X115 flash_0.x7.dcgint.t10 flash_0.x7.pos_en_b.t6 VGND.t42 VGND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X116 a_20416_28577# flash_0.x7.neg_mid_b.t10 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X117 flash_0.x7.VOUT.t11 flash_0.x7.neg_mid_b.t11 flash_0.x7.dcgint.t5 flash_0.x7.dcgint.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X118 VDPWR.t17 ui_in[0].t14 flash_0.x7.neg_mid VDPWR.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X119 flash_0.x7.neg_mid_b.t1 flash_0.x7.neg_en_b.t8 VDPWR.t55 VDPWR.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X120 flash_0.x4.neg_en_b.t1 ui_in[1].t14 VGND.t16 VGND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X121 flash_0.x4.pos_en_b.t2 ui_in[0].t15 VGND.t3 VGND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X122 flash_0.x4.neg_mid ui_in[1].t15 VDPWR.t26 VDPWR.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X123 VDPWR.t1 ui_in[0].t16 flash_0.x7.neg_en_b.t0 VDPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X124 flash_0.x7.dcgint.t4 flash_0.x7.neg_mid_b.t12 flash_0.x7.VOUT.t12 flash_0.x7.dcgint.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X125 flash_0.x2.clkinb clk.t3 VGND.t21 VGND.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X126 flash_0.x7.VOUT.t13 flash_0.x7.neg_mid_b.t13 flash_0.x7.dcgint.t3 flash_0.x7.dcgint.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X127 flash_0.x4.VOUT.t3 VDPWR.t69 flash_0.x4.vintp flash_0.x7.VPRGPOS.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X128 flash_0.x7.dcgint.t9 flash_0.x7.pos_en_b.t6 VGND.t40 VGND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X129 flash_0.x3.clka.t1 flash_0.x3.clkina VGND.t46 VGND.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X130 flash_0.x5.A.t2 flash_0.x5.A.t0 a_9352_28387# flash_0.x5.A.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.5
X131 flash_0.x7.dcgint.t1 flash_0.x7.neg_mid_b.t14 flash_0.x7.VOUT.t10 flash_0.x7.dcgint.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X132 flash_0.x7.neg_mid_b.t0 flash_0.x7.neg_en_b.t9 VDPWR.t15 VDPWR.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X133 flash_0.x7.vintp VDPWR.t70 flash_0.x7.VOUT.t6 flash_0.x7.VPRGPOS.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X134 flash_0.x4.neg_en_b.t0 ui_in[1].t16 VDPWR.t24 VDPWR.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=3
X135 flash_0.x4.pos_en_b.t0 ui_in[0].t17 VDPWR.t11 VDPWR.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X136 VGND.t8 flash_0.x4.pos_en_b.t6 flash_0.x4.pos_mid VGND.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X137 flash_0.x7.VPRGNEG flash_0.x7.neg_mid_b.t15 flash_0.x7.neg_mid flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.145 ps=1.58 w=0.5 l=1
X138 flash_0.x7.VOUT.t5 VDPWR.t71 flash_0.x7.vintp flash_0.x7.VPRGPOS.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X139 flash_0.x2.stage2 flash_0.x2.stage2 flash_0.x2.stage1 flash_0.x2.stage2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X140 flash_0.x7.VPRGPOS.t30 flash_0.x4.pos_mid_b.t8 flash_0.x4.vintp flash_0.x7.VPRGPOS.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X141 flash_0.x4.neg_mid ui_in[1].t17 VDPWR.t22 VDPWR.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X142 flash_0.x7.vintp flash_0.x7.pos_mid_b.t7 flash_0.x7.VPRGPOS.t20 flash_0.x7.VPRGPOS.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X143 flash_0.x7.VOUT.t4 VDPWR.t72 flash_0.x7.vintp flash_0.x7.VPRGPOS.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X144 flash_0.x7.VPRGPOS.t19 flash_0.x7.pos_mid_b flash_0.x7.pos_mid flash_0.x7.VPRGPOS.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X145 flash_0.x7.VPRGPOS.t27 flash_0.x4.pos_mid_b flash_0.x4.pos_mid flash_0.x7.VPRGPOS.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X146 VGND.t7 flash_0.x4.pos_en_b.t6 flash_0.x4.pos_mid VGND.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X147 uo_out[0].t1 flash_0.x5.A.t5 VGND.t26 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X148 flash_0.x3.clkina flash_0.x3.clkinb VGND.t57 VGND.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X149 flash_0.x7.vintp VDPWR.t73 flash_0.x7.VOUT.t3 flash_0.x7.VPRGPOS.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X150 flash_0.x7.VPRGPOS.t17 flash_0.x7.pos_mid_b.t8 flash_0.x7.vintp flash_0.x7.VPRGPOS.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X151 flash_0.x6.Y ui_in[2].t2 VDPWR.t13 VDPWR.t12 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X152 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG flash_0.x2.stage2 flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
R0 VGND.t28 VGND.n108 1.77808e+07
R1 VGND.n211 VGND.n210 1.32662e+07
R2 VGND.n108 VGND.t39 9.06413e+06
R3 VGND.n211 VGND.n24 7.77048e+06
R4 VGND.n126 VGND.n116 136400
R5 VGND.n123 VGND.n98 77206.1
R6 VGND.n178 VGND.n63 55379.3
R7 VGND.n128 VGND.n127 41452.9
R8 VGND.n124 VGND.n122 28158.7
R9 VGND.n82 VGND.n67 26564
R10 VGND.n131 VGND.n116 26182
R11 VGND.n82 VGND.n81 19464
R12 VGND.n127 VGND.n126 18707.2
R13 VGND.n177 VGND.n176 17794
R14 VGND.n212 VGND.n22 17579
R15 VGND.n45 VGND.n41 17010.2
R16 VGND.n52 VGND.n41 17010.2
R17 VGND.n189 VGND.n56 17010.2
R18 VGND.n180 VGND.n56 17010.2
R19 VGND.n150 VGND.n116 16052.9
R20 VGND.n124 VGND.n22 15944.1
R21 VGND.n176 VGND.n82 15655.2
R22 VGND.n123 VGND.n99 15267.5
R23 VGND.n178 VGND.n177 13983.9
R24 VGND.n177 VGND.n64 12678.4
R25 VGND.n126 VGND.n125 11203.8
R26 VGND.n213 VGND.n212 8682.25
R27 VGND.n153 VGND.n99 8288.46
R28 VGND.n71 VGND.n22 7672.91
R29 VGND.n115 VGND.t32 6465.71
R30 VGND.n125 VGND.n123 5878.85
R31 VGND.n211 VGND.n23 5801.34
R32 VGND.n58 VGND.n55 5607.68
R33 VGND.n43 VGND.n40 5607.68
R34 VGND.n40 VGND.n23 5607.68
R35 VGND.n62 VGND.n55 5607.68
R36 VGND.n101 VGND.n100 5067.26
R37 VGND.n129 VGND.n128 4557.14
R38 VGND.t36 VGND.t22 4288.33
R39 VGND.t22 VGND.t17 4288.33
R40 VGND.t6 VGND.t2 4288.33
R41 VGND.t2 VGND.t4 4288.33
R42 VGND.n174 VGND.n83 3957.38
R43 VGND.n174 VGND.n84 3957.38
R44 VGND.n120 VGND.n84 3957.38
R45 VGND.n120 VGND.n83 3957.38
R46 VGND.n72 VGND.n68 3957.38
R47 VGND.n72 VGND.n69 3957.38
R48 VGND.n80 VGND.n69 3957.38
R49 VGND.n80 VGND.n68 3957.38
R50 VGND.n209 VGND.n25 3790.36
R51 VGND.n60 VGND.n25 3790.36
R52 VGND.n195 VGND.n194 3790.36
R53 VGND.n194 VGND.n38 3790.36
R54 VGND.t0 VGND.n152 3495.43
R55 VGND.n130 VGND.t12 3495.43
R56 VGND.n81 VGND.t14 3200.66
R57 VGND.n71 VGND.t14 3200.66
R58 VGND.n152 VGND.n98 2827
R59 VGND.n131 VGND.n130 2827
R60 VGND.n43 VGND.n39 2736.73
R61 VGND.n151 VGND.n150 2648.22
R62 VGND.n127 VGND.n122 2546
R63 VGND.t17 VGND.n151 2345.18
R64 VGND.t4 VGND.n129 2345.18
R65 VGND.n178 VGND.n62 2341.85
R66 VGND.n153 VGND.t0 2331.85
R67 VGND.n63 VGND.n58 2309.11
R68 VGND.n54 VGND.n53 2233.78
R69 VGND.n125 VGND.n124 2176.84
R70 VGND.n212 VGND.n211 1977.24
R71 VGND.n214 VGND.n20 1900.12
R72 VGND.n214 VGND.n21 1900.12
R73 VGND.n66 VGND.n21 1900.12
R74 VGND.n66 VGND.n20 1900.12
R75 VGND.n191 VGND.n190 1830.35
R76 VGND.t12 VGND.n115 1820.3
R77 VGND.n128 VGND.n64 1788.04
R78 VGND.n122 VGND.n121 1768.36
R79 VGND.n44 VGND.n23 1501.04
R80 VGND.n54 VGND.n39 1195.35
R81 VGND.n176 VGND.n175 1151.51
R82 VGND.n51 VGND.n42 1139.95
R83 VGND.n46 VGND.n42 1139.95
R84 VGND.n188 VGND.n57 1139.95
R85 VGND.n181 VGND.n57 1139.95
R86 VGND.t43 VGND.n99 1094.37
R87 VGND.n121 VGND.t25 1089.55
R88 VGND.n175 VGND.t25 1089.55
R89 VGND.n101 VGND.n54 931.699
R90 VGND.n62 VGND.n61 883.615
R91 VGND.n152 VGND.t36 792.894
R92 VGND.n130 VGND.t6 792.894
R93 VGND.t52 VGND.t62 757.616
R94 VGND.n67 VGND.t66 660
R95 VGND.n213 VGND.t66 660
R96 VGND.n179 VGND.n58 657.409
R97 VGND.n15 VGND.t50 650.87
R98 VGND.t54 VGND.t20 597.753
R99 VGND.n149 VGND.n132 535.718
R100 VGND.n155 VGND.n154 535.718
R101 VGND.n108 VGND.n101 522.082
R102 VGND.t32 VGND.t30 487.856
R103 VGND.n61 VGND.t52 478.974
R104 VGND.t45 VGND.t58 470.42
R105 VGND.n208 VGND.n207 437.836
R106 VGND.n207 VGND.n27 437.836
R107 VGND.n197 VGND.n37 437.836
R108 VGND.n197 VGND.n196 437.836
R109 VGND.n210 VGND.t20 424.973
R110 VGND.n44 VGND.n43 417.728
R111 VGND.n191 VGND.n54 402.44
R112 VGND.t62 VGND.n59 378.808
R113 VGND.n59 VGND.t54 378.808
R114 VGND.t56 VGND.t10 350.719
R115 VGND.n114 VGND.t28 304.329
R116 VGND.t58 VGND.n192 297.404
R117 VGND.n119 VGND.n118 257.13
R118 VGND.n119 VGND.n86 257.13
R119 VGND.n79 VGND.n70 257.13
R120 VGND.n79 VGND.n78 257.13
R121 VGND.n193 VGND.t45 235.209
R122 VGND.n112 VGND.t29 230.898
R123 VGND.n109 VGND.t31 230.898
R124 VGND.n110 VGND.t33 230.898
R125 VGND.n105 VGND.t40 230.898
R126 VGND.n102 VGND.t42 230.898
R127 VGND.n103 VGND.t44 230.898
R128 VGND.n118 VGND.n85 229.272
R129 VGND.n172 VGND.n86 229.272
R130 VGND.n74 VGND.n70 229.272
R131 VGND.n78 VGND.n77 229.272
R132 VGND.n199 VGND.t57 227.643
R133 VGND.n205 VGND.t55 227.643
R134 VGND.n26 VGND.t21 227.398
R135 VGND.n34 VGND.t11 227.398
R136 VGND.n193 VGND.t56 222.901
R137 VGND.n215 VGND.n19 221.742
R138 VGND.n65 VGND.n19 221.742
R139 VGND.n65 VGND.n18 221.742
R140 VGND.t10 VGND.n24 221.728
R141 VGND.n132 VGND.n131 188.038
R142 VGND.n155 VGND.n98 188.038
R143 VGND.t30 VGND.n114 183.528
R144 VGND.n150 VGND.n149 180.132
R145 VGND.n154 VGND.n153 180.132
R146 VGND.t41 VGND.t43 157.787
R147 VGND.n216 VGND.n18 152.194
R148 VGND.n151 VGND.n90 152.111
R149 VGND.n129 VGND.n117 152.111
R150 VGND.n122 VGND.n64 147.569
R151 VGND.n20 VGND.n18 146.25
R152 VGND.t66 VGND.n20 146.25
R153 VGND.n21 VGND.n19 146.25
R154 VGND.t66 VGND.n21 146.25
R155 VGND.n120 VGND.n119 117.001
R156 VGND.n121 VGND.n120 117.001
R157 VGND.n174 VGND.n173 117.001
R158 VGND.n175 VGND.n174 117.001
R159 VGND.n80 VGND.n79 117.001
R160 VGND.n81 VGND.n80 117.001
R161 VGND.n73 VGND.n72 117.001
R162 VGND.n72 VGND.n71 117.001
R163 VGND.n192 VGND.n191 107.427
R164 VGND.n53 VGND.n40 102.35
R165 VGND.n190 VGND.n55 102.35
R166 VGND.t39 VGND.n107 98.4295
R167 VGND.n60 VGND.n27 97.5005
R168 VGND.n61 VGND.n60 97.5005
R169 VGND.n209 VGND.n208 97.5005
R170 VGND.n210 VGND.n209 97.5005
R171 VGND.n38 VGND.n37 97.5005
R172 VGND.n192 VGND.n38 97.5005
R173 VGND.n196 VGND.n195 97.5005
R174 VGND.n195 VGND.n24 97.5005
R175 VGND.n163 VGND.n162 97.1505
R176 VGND.n96 VGND.n95 97.1505
R177 VGND.n159 VGND.n158 97.1505
R178 VGND.n92 VGND.n91 97.1505
R179 VGND.n161 VGND.n160 97.1505
R180 VGND.n94 VGND.n93 97.1505
R181 VGND.n145 VGND.n144 97.1505
R182 VGND.n138 VGND.n137 97.1505
R183 VGND.n141 VGND.n140 97.1505
R184 VGND.n134 VGND.n133 97.1505
R185 VGND.n143 VGND.n142 97.1505
R186 VGND.n136 VGND.n135 97.1505
R187 VGND.n100 VGND.n63 95.855
R188 VGND.n162 VGND.t47 95.7605
R189 VGND.n162 VGND.t34 95.7605
R190 VGND.n95 VGND.t1 95.7605
R191 VGND.n95 VGND.t70 95.7605
R192 VGND.n158 VGND.t23 95.7605
R193 VGND.n158 VGND.t60 95.7605
R194 VGND.n91 VGND.t35 95.7605
R195 VGND.n91 VGND.t37 95.7605
R196 VGND.n160 VGND.t24 95.7605
R197 VGND.n160 VGND.t18 95.7605
R198 VGND.n93 VGND.t61 95.7605
R199 VGND.n93 VGND.t38 95.7605
R200 VGND.n144 VGND.t3 95.7605
R201 VGND.n144 VGND.t48 95.7605
R202 VGND.n137 VGND.t16 95.7605
R203 VGND.n137 VGND.t9 95.7605
R204 VGND.n140 VGND.t64 95.7605
R205 VGND.n140 VGND.t68 95.7605
R206 VGND.n133 VGND.t27 95.7605
R207 VGND.n133 VGND.t7 95.7605
R208 VGND.n142 VGND.t65 95.7605
R209 VGND.n142 VGND.t5 95.7605
R210 VGND.n135 VGND.t13 95.7605
R211 VGND.n135 VGND.t8 95.7605
R212 VGND.n170 VGND.t26 83.754
R213 VGND.n76 VGND.t15 83.7172
R214 VGND.n36 VGND.t59 83.1807
R215 VGND.n28 VGND.t53 83.1807
R216 VGND.n35 VGND.t46 82.9558
R217 VGND.n29 VGND.t63 82.9558
R218 VGND.n30 VGND.t19 82.8472
R219 VGND.n107 VGND.n106 73.7068
R220 VGND.n114 VGND.n113 73.7068
R221 VGND.n66 VGND.n65 65.0005
R222 VGND.n67 VGND.n66 65.0005
R223 VGND.n215 VGND.n214 65.0005
R224 VGND.n214 VGND.n213 65.0005
R225 VGND.n107 VGND.t41 59.3584
R226 VGND.n216 VGND.n215 56.9466
R227 VGND.n118 VGND.n83 53.1823
R228 VGND.n83 VGND.t25 53.1823
R229 VGND.n86 VGND.n84 53.1823
R230 VGND.n84 VGND.t25 53.1823
R231 VGND.n70 VGND.n68 53.1823
R232 VGND.n68 VGND.t14 53.1823
R233 VGND.n78 VGND.n69 53.1823
R234 VGND.n69 VGND.t14 53.1823
R235 VGND.n217 VGND.t67 41.2645
R236 VGND.n173 VGND.n85 27.8593
R237 VGND.n173 VGND.n172 27.8593
R238 VGND.n74 VGND.n73 27.8593
R239 VGND.n77 VGND.n73 27.8593
R240 VGND.n57 VGND.n56 26.5914
R241 VGND.n100 VGND.n56 26.5914
R242 VGND.n42 VGND.n41 26.5914
R243 VGND.n41 VGND.n39 26.5914
R244 VGND.n207 VGND.n25 24.3755
R245 VGND.n59 VGND.n25 24.3755
R246 VGND.n197 VGND.n194 24.3755
R247 VGND.n194 VGND.n193 24.3755
R248 VGND.n179 VGND.n178 20.4593
R249 VGND.n75 VGND.n74 9.35514
R250 VGND.n77 VGND 9.33194
R251 VGND.n172 VGND.n171 9.3005
R252 VGND.n171 VGND.n85 9.3005
R253 VGND.n46 VGND.n45 9.28621
R254 VGND.n45 VGND.n44 9.28621
R255 VGND.n189 VGND.n188 9.28621
R256 VGND.n190 VGND.n189 9.28621
R257 VGND.n52 VGND.n51 9.28621
R258 VGND.n53 VGND.n52 9.28621
R259 VGND.n181 VGND.n180 9.28621
R260 VGND.n180 VGND.n179 9.28621
R261 VGND.n219 VGND.n16 8.39735
R262 VGND.n48 VGND.n47 8.21246
R263 VGND.n187 VGND.n186 8.21246
R264 VGND.n49 VGND.n48 7.33652
R265 VGND.n186 VGND.n185 7.33652
R266 VGND.n165 VGND.n90 6.24424
R267 VGND.n117 VGND.n87 6.24424
R268 VGND.n148 VGND.n147 6.00831
R269 VGND.n157 VGND.n156 5.96627
R270 VGND.n47 VGND 5.82387
R271 VGND.n187 VGND 5.82387
R272 VGND.n218 VGND.n217 5.18907
R273 VGND.n50 VGND 5.15194
R274 VGND.n182 VGND 5.15194
R275 VGND.n170 VGND.n169 5.15155
R276 VGND.n15 VGND.t49 4.756
R277 VGND.n111 VGND.n110 4.5005
R278 VGND.n111 VGND.n109 4.5005
R279 VGND.n112 VGND.n111 4.5005
R280 VGND.n104 VGND.n103 4.5005
R281 VGND.n104 VGND.n102 4.5005
R282 VGND.n105 VGND.n104 4.5005
R283 VGND.n33 VGND.n32 4.12801
R284 VGND.n184 VGND.n183 4.12801
R285 VGND.n151 VGND.n115 4.11265
R286 VGND.n202 VGND 3.81988
R287 VGND.n221 VGND 3.32011
R288 VGND.n37 VGND.n36 3.31952
R289 VGND.n28 VGND.n27 3.31952
R290 VGND.n201 VGND.n33 3.218
R291 VGND.n16 VGND.n15 3.20171
R292 VGND.n166 VGND.n89 3.12737
R293 VGND.n168 VGND.n167 3.00925
R294 VGND.n156 VGND.n155 2.81159
R295 VGND.n148 VGND.n132 2.79528
R296 uio_oe[7] VGND.n221 2.60868
R297 VGND VGND.n148 2.41626
R298 VGND.n156 VGND 2.39996
R299 VGND.n149 VGND 2.3442
R300 VGND.n154 VGND 2.3442
R301 VGND.n217 VGND.n216 2.3255
R302 VGND.n139 VGND.n136 2.2505
R303 VGND.n146 VGND.n143 2.2505
R304 VGND.n139 VGND.n134 2.2505
R305 VGND.n146 VGND.n141 2.2505
R306 VGND.n139 VGND.n138 2.2505
R307 VGND.n146 VGND.n145 2.2505
R308 VGND.n97 VGND.n94 2.2505
R309 VGND.n164 VGND.n161 2.2505
R310 VGND.n97 VGND.n92 2.2505
R311 VGND.n164 VGND.n159 2.2505
R312 VGND.n97 VGND.n96 2.2505
R313 VGND.n164 VGND.n163 2.2505
R314 VGND.n113 VGND.n112 2.04916
R315 VGND.n106 VGND.n105 2.04916
R316 VGND.n169 VGND.n168 2.00487
R317 VGND.n184 VGND.n31 1.913
R318 VGND.n169 VGND.n17 1.74613
R319 VGND.n31 VGND.n30 1.5555
R320 VGND.n208 VGND.n26 1.5505
R321 VGND.n196 VGND.n34 1.5505
R322 VGND.n166 VGND.n165 1.31425
R323 VGND.n203 VGND.n31 1.3055
R324 VGND.n168 VGND.n87 1.248
R325 VGND.n218 VGND.n17 1.188
R326 VGND.n202 VGND.n17 1.1555
R327 VGND.n36 VGND.n35 0.879043
R328 VGND.n29 VGND.n28 0.879043
R329 VGND.n221 VGND.n220 0.751794
R330 VGND.n219 VGND.n218 0.525188
R331 VGND.n204 VGND.n203 0.501003
R332 VGND.n201 VGND.n200 0.501003
R333 VGND.n48 VGND.n42 0.443357
R334 VGND.n186 VGND.n57 0.443357
R335 VGND.n207 VGND.n206 0.404848
R336 VGND.n198 VGND.n197 0.404848
R337 VGND.n164 VGND.n157 0.36615
R338 VGND.n147 VGND.n146 0.365657
R339 VGND.n106 VGND.n89 0.285933
R340 VGND.n113 VGND.n88 0.28175
R341 VGND.n167 VGND.n166 0.27425
R342 VGND.n167 VGND.n88 0.236484
R343 VGND.n206 VGND.n205 0.221088
R344 VGND.n199 VGND.n198 0.221088
R345 VGND.n205 VGND 0.214961
R346 VGND VGND.n199 0.214961
R347 VGND.n111 VGND 0.204732
R348 VGND.n104 VGND 0.204732
R349 VGND VGND.n202 0.177375
R350 VGND.n75 VGND.n16 0.168469
R351 VGND.n220 VGND.n219 0.166437
R352 VGND.n0 uo_out[1] 0.16627
R353 VGND.n1 uo_out[2] 0.16627
R354 VGND.n2 uo_out[3] 0.16627
R355 VGND.n3 uo_out[4] 0.16627
R356 VGND.n4 uo_out[5] 0.16627
R357 VGND.n5 uo_out[6] 0.16627
R358 VGND.n6 uo_out[7] 0.16627
R359 VGND.n7 uio_out[0] 0.16627
R360 VGND.n8 uio_out[1] 0.16627
R361 VGND.n9 uio_out[2] 0.16627
R362 VGND.n10 uio_out[3] 0.16627
R363 VGND.n11 uio_out[4] 0.16627
R364 VGND.n12 uio_out[5] 0.16627
R365 VGND.n13 uio_out[6] 0.16627
R366 VGND.n14 uio_out[7] 0.16627
R367 uio_oe[0] VGND.n228 0.16627
R368 uio_oe[1] VGND.n227 0.16627
R369 uio_oe[2] VGND.n226 0.16627
R370 uio_oe[3] VGND.n225 0.16627
R371 uio_oe[4] VGND.n224 0.16627
R372 uio_oe[5] VGND.n223 0.16627
R373 uio_oe[6] VGND.n222 0.16627
R374 VGND.n90 VGND 0.157483
R375 VGND.n117 VGND 0.157483
R376 VGND.n50 VGND.n49 0.15675
R377 VGND.n185 VGND.n182 0.15675
R378 VGND.n47 VGND.n46 0.1555
R379 VGND.n51 VGND.n50 0.1555
R380 VGND.n188 VGND.n187 0.1555
R381 VGND.n182 VGND.n181 0.1555
R382 VGND.n163 VGND 0.102773
R383 VGND.n96 VGND 0.102773
R384 VGND.n159 VGND 0.102773
R385 VGND.n92 VGND 0.102773
R386 VGND.n161 VGND 0.102773
R387 VGND.n94 VGND 0.102773
R388 VGND.n145 VGND 0.102773
R389 VGND.n138 VGND 0.102773
R390 VGND.n141 VGND 0.102773
R391 VGND.n134 VGND 0.102773
R392 VGND.n143 VGND 0.102773
R393 VGND.n136 VGND 0.102773
R394 VGND.n204 VGND.n26 0.0904491
R395 VGND.n200 VGND.n34 0.0904491
R396 VGND VGND.n204 0.0659475
R397 VGND.n200 VGND 0.0659475
R398 VGND.n49 VGND.n33 0.0657174
R399 VGND.n185 VGND.n184 0.0657174
R400 VGND.n220 VGND 0.062375
R401 VGND.n30 VGND 0.0609396
R402 VGND VGND.n201 0.05925
R403 VGND.n203 VGND 0.05925
R404 VGND.n109 VGND 0.0544773
R405 VGND.n110 VGND 0.0544773
R406 VGND.n102 VGND 0.0544773
R407 VGND.n103 VGND 0.0544773
R408 VGND.n112 VGND 0.048
R409 VGND.n105 VGND 0.048
R410 VGND.n171 VGND.n170 0.034875
R411 VGND.n183 VGND.t51 0.0314016
R412 VGND.n32 VGND.t69 0.0314016
R413 VGND VGND.n88 0.0312579
R414 VGND.n0 uo_out[2] 0.0302667
R415 VGND.n1 uo_out[3] 0.0302667
R416 VGND.n2 uo_out[4] 0.0302667
R417 VGND.n3 uo_out[5] 0.0302667
R418 VGND.n4 uo_out[6] 0.0302667
R419 VGND.n5 uo_out[7] 0.0302667
R420 VGND.n6 uio_out[0] 0.0302667
R421 VGND.n7 uio_out[1] 0.0302667
R422 VGND.n8 uio_out[2] 0.0302667
R423 VGND.n9 uio_out[3] 0.0302667
R424 VGND.n10 uio_out[4] 0.0302667
R425 VGND.n11 uio_out[5] 0.0302667
R426 VGND.n12 uio_out[6] 0.0302667
R427 VGND.n13 uio_out[7] 0.0302667
R428 VGND.n14 uio_oe[0] 0.0302667
R429 VGND.n228 uio_oe[1] 0.0302667
R430 VGND.n227 uio_oe[2] 0.0302667
R431 VGND.n226 uio_oe[3] 0.0302667
R432 VGND.n225 uio_oe[4] 0.0302667
R433 VGND.n224 uio_oe[5] 0.0302667
R434 VGND.n223 uio_oe[6] 0.0302667
R435 VGND.n222 uio_oe[7] 0.0302667
R436 VGND VGND.n89 0.0270748
R437 VGND VGND.n76 0.0244521
R438 VGND.n206 VGND.n29 0.0194951
R439 VGND.n198 VGND.n35 0.0194951
R440 VGND.n146 VGND.n87 0.0182165
R441 VGND.n165 VGND.n164 0.0182165
R442 VGND.n147 VGND.n139 0.0132953
R443 VGND.n157 VGND.n97 0.0128031
R444 uo_out[2] VGND.n0 0.010027
R445 uo_out[3] VGND.n1 0.010027
R446 uo_out[4] VGND.n2 0.010027
R447 uo_out[5] VGND.n3 0.010027
R448 uo_out[6] VGND.n4 0.010027
R449 uo_out[7] VGND.n5 0.010027
R450 uio_out[0] VGND.n6 0.010027
R451 uio_out[1] VGND.n7 0.010027
R452 uio_out[2] VGND.n8 0.010027
R453 uio_out[3] VGND.n9 0.010027
R454 uio_out[4] VGND.n10 0.010027
R455 uio_out[5] VGND.n11 0.010027
R456 uio_out[6] VGND.n12 0.010027
R457 uio_out[7] VGND.n13 0.010027
R458 uio_oe[0] VGND.n14 0.010027
R459 VGND.n228 uio_oe[1] 0.010027
R460 VGND.n227 uio_oe[2] 0.010027
R461 VGND.n226 uio_oe[3] 0.010027
R462 VGND.n225 uio_oe[4] 0.010027
R463 VGND.n224 uio_oe[5] 0.010027
R464 VGND.n223 uio_oe[6] 0.010027
R465 VGND.n222 uio_oe[7] 0.010027
R466 VGND.n171 VGND 0.008625
R467 VGND.n76 VGND.n75 0.0012485
R468 VGND.n183 VGND 0.000981102
R469 VGND.n32 VGND 0.000981102
R470 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t1 649.691
R471 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t0 227.442
R472 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t2 227.361
R473 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t7 216.731
R474 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t8 216.731
R475 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t6 216.731
R476 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t3 216.731
R477 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t4 216.731
R478 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t5 216.731
R479 flash_0.x7.VPRGPOS.n6 flash_0.x7.VPRGPOS.n4 4689.72
R480 flash_0.x7.VPRGPOS.n9 flash_0.x7.VPRGPOS.n8 4689.72
R481 flash_0.x7.VPRGPOS.n7 flash_0.x7.VPRGPOS.n6 1828.1
R482 flash_0.x7.VPRGPOS.n9 flash_0.x7.VPRGPOS.n3 1828.1
R483 flash_0.x7.VPRGPOS.n5 flash_0.x7.VPRGPOS.n1 902.777
R484 flash_0.x7.VPRGPOS.n5 flash_0.x7.VPRGPOS.n2 902.777
R485 flash_0.x7.VPRGPOS.n10 flash_0.x7.VPRGPOS.n2 880.232
R486 flash_0.x7.VPRGPOS.n11 flash_0.x7.VPRGPOS.n1 874.658
R487 flash_0.x7.VPRGPOS.t0 flash_0.x7.VPRGPOS.t18 809.375
R488 flash_0.x7.VPRGPOS.t2 flash_0.x7.VPRGPOS.t6 809.375
R489 flash_0.x7.VPRGPOS.n12 flash_0.x7.VPRGPOS.t29 649.856
R490 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t30 649.715
R491 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t22 649.715
R492 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t26 649.691
R493 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t19 649.691
R494 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t7 649.691
R495 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t27 649.691
R496 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t5 649.691
R497 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t20 649.691
R498 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n14 594.301
R499 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n13 594.301
R500 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n18 594.301
R501 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n19 594.301
R502 flash_0.x7.VPRGPOS.t8 flash_0.x7.VPRGPOS.t12 246.875
R503 flash_0.x7.VPRGPOS.t24 flash_0.x7.VPRGPOS.t8 246.875
R504 flash_0.x7.VPRGPOS.t14 flash_0.x7.VPRGPOS.t24 246.875
R505 flash_0.x7.VPRGPOS.t1 flash_0.x7.VPRGPOS.t14 246.875
R506 flash_0.x7.VPRGPOS.t15 flash_0.x7.VPRGPOS.t13 246.875
R507 flash_0.x7.VPRGPOS.t3 flash_0.x7.VPRGPOS.t15 246.875
R508 flash_0.x7.VPRGPOS.t9 flash_0.x7.VPRGPOS.t3 246.875
R509 flash_0.x7.VPRGPOS.t31 flash_0.x7.VPRGPOS.t9 246.875
R510 flash_0.x7.VPRGPOS.n0 flash_0.x7.VPRGPOS.t1 237.5
R511 flash_0.x7.VPRGPOS.n15 flash_0.x7.VPRGPOS.t31 237.5
R512 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t11 82.8472
R513 flash_0.x7.VPRGPOS.n14 flash_0.x7.VPRGPOS.t10 55.3905
R514 flash_0.x7.VPRGPOS.n14 flash_0.x7.VPRGPOS.t32 55.3905
R515 flash_0.x7.VPRGPOS.n13 flash_0.x7.VPRGPOS.t16 55.3905
R516 flash_0.x7.VPRGPOS.n13 flash_0.x7.VPRGPOS.t4 55.3905
R517 flash_0.x7.VPRGPOS.n18 flash_0.x7.VPRGPOS.t21 55.3905
R518 flash_0.x7.VPRGPOS.n18 flash_0.x7.VPRGPOS.t17 55.3905
R519 flash_0.x7.VPRGPOS.n19 flash_0.x7.VPRGPOS.t23 55.3905
R520 flash_0.x7.VPRGPOS.n19 flash_0.x7.VPRGPOS.t25 55.3905
R521 flash_0.x7.VPRGPOS.n6 flash_0.x7.VPRGPOS.n5 37.0005
R522 flash_0.x7.VPRGPOS.n10 flash_0.x7.VPRGPOS.n9 37.0005
R523 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n0 16.1367
R524 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n15 16.1367
R525 flash_0.x7.VPRGPOS.n17 flash_0.x7.VPRGPOS 13.9898
R526 flash_0.x7.VPRGPOS.n0 flash_0.x7.VPRGPOS.t0 9.3755
R527 flash_0.x7.VPRGPOS.n15 flash_0.x7.VPRGPOS.t2 9.3755
R528 flash_0.x7.VPRGPOS.n4 flash_0.x7.VPRGPOS.n1 3.03329
R529 flash_0.x7.VPRGPOS.n8 flash_0.x7.VPRGPOS.n2 3.03329
R530 flash_0.x7.VPRGPOS.n16 flash_0.x7.VPRGPOS 2.77904
R531 flash_0.x7.VPRGPOS.n11 flash_0.x7.VPRGPOS.n10 2.70819
R532 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n17 2.54902
R533 flash_0.x7.VPRGPOS.n12 flash_0.x7.VPRGPOS.n11 1.8605
R534 flash_0.x7.VPRGPOS.n4 flash_0.x7.VPRGPOS.n3 1.85038
R535 flash_0.x7.VPRGPOS.n8 flash_0.x7.VPRGPOS.n7 1.85038
R536 flash_0.x7.VPRGPOS.n16 flash_0.x7.VPRGPOS.n12 1.79707
R537 flash_0.x7.VPRGPOS.n17 flash_0.x7.VPRGPOS.n16 1.40849
R538 flash_0.x7.VPRGPOS.t28 flash_0.x7.VPRGPOS.n3 1.18321
R539 flash_0.x7.VPRGPOS.n7 flash_0.x7.VPRGPOS.t28 1.18321
R540 VAPWR.n62 VAPWR.n4 2380.24
R541 VAPWR.n114 VAPWR.n73 2380.24
R542 VAPWR.n64 VAPWR.n4 2376.31
R543 VAPWR.n116 VAPWR.n73 2376.31
R544 VAPWR.n44 VAPWR.n42 2332.91
R545 VAPWR.n45 VAPWR.n44 2332.91
R546 VAPWR.n46 VAPWR.n45 2332.91
R547 VAPWR.n46 VAPWR.n42 2332.91
R548 VAPWR.n27 VAPWR.n25 2332.91
R549 VAPWR.n28 VAPWR.n27 2332.91
R550 VAPWR.n29 VAPWR.n28 2332.91
R551 VAPWR.n29 VAPWR.n25 2332.91
R552 VAPWR.n13 VAPWR.n12 2332.91
R553 VAPWR.n13 VAPWR.n11 2332.91
R554 VAPWR.n93 VAPWR.n92 2332.91
R555 VAPWR.n93 VAPWR.n91 2332.91
R556 VAPWR.n87 VAPWR.n83 1577.4
R557 VAPWR.n84 VAPWR.n81 1577.4
R558 VAPWR.n47 VAPWR.n38 1551.32
R559 VAPWR.n43 VAPWR.n38 1551.32
R560 VAPWR.n26 VAPWR.n24 1551.32
R561 VAPWR.n26 VAPWR.n21 1551.32
R562 VAPWR.n30 VAPWR.n21 1551.32
R563 VAPWR.n30 VAPWR.n24 1551.32
R564 VAPWR.n47 VAPWR.n41 1538.26
R565 VAPWR.n43 VAPWR.n41 1538.26
R566 VAPWR.n58 VAPWR.n7 1516.38
R567 VAPWR.n58 VAPWR.n6 1516.38
R568 VAPWR.n110 VAPWR.n76 1516.38
R569 VAPWR.n110 VAPWR.n75 1516.38
R570 VAPWR.n14 VAPWR.n7 1514.88
R571 VAPWR.n14 VAPWR.n6 1514.88
R572 VAPWR.n94 VAPWR.n76 1514.88
R573 VAPWR.n94 VAPWR.n75 1514.88
R574 VAPWR.n12 VAPWR.n5 1046.2
R575 VAPWR.n11 VAPWR.n5 1046.2
R576 VAPWR.n92 VAPWR.n74 1046.2
R577 VAPWR.n91 VAPWR.n74 1046.2
R578 VAPWR.n85 VAPWR.n84 722.497
R579 VAPWR.n87 VAPWR.n86 722.497
R580 VAPWR.n0 VAPWR.t10 649.99
R581 VAPWR.n121 VAPWR.t14 649.99
R582 VAPWR.n1 VAPWR.t6 649.765
R583 VAPWR.n71 VAPWR.t1 649.765
R584 VAPWR.t5 VAPWR.t9 487.901
R585 VAPWR.t0 VAPWR.t13 487.901
R586 VAPWR.n66 VAPWR.n3 460.425
R587 VAPWR.n118 VAPWR.n72 460.425
R588 VAPWR.n66 VAPWR.n65 459.671
R589 VAPWR.n118 VAPWR.n117 459.671
R590 VAPWR.n40 VAPWR.n37 386.635
R591 VAPWR.n48 VAPWR.n40 386.635
R592 VAPWR.n49 VAPWR.n37 386.635
R593 VAPWR.n23 VAPWR.n20 386.635
R594 VAPWR.n31 VAPWR.n23 386.635
R595 VAPWR.n32 VAPWR.n20 386.635
R596 VAPWR.n15 VAPWR.n8 386.635
R597 VAPWR.n15 VAPWR.n9 386.635
R598 VAPWR.n57 VAPWR.n8 386.635
R599 VAPWR.n57 VAPWR.n9 386.635
R600 VAPWR.n95 VAPWR.n77 386.635
R601 VAPWR.n95 VAPWR.n78 386.635
R602 VAPWR.n109 VAPWR.n78 386.635
R603 VAPWR.n109 VAPWR.n77 386.635
R604 VAPWR.n64 VAPWR.t5 331.582
R605 VAPWR.n116 VAPWR.t0 331.582
R606 VAPWR.n61 VAPWR.n60 251.28
R607 VAPWR.n113 VAPWR.n112 251.28
R608 VAPWR.t2 VAPWR 236.188
R609 VAPWR.n97 VAPWR.t2 236.011
R610 VAPWR.n49 VAPWR 195.012
R611 VAPWR.n32 VAPWR 195.012
R612 VAPWR VAPWR.n48 191.625
R613 VAPWR VAPWR.n31 191.625
R614 VAPWR.n106 VAPWR.n82 184.847
R615 VAPWR.n107 VAPWR.n106 184.847
R616 VAPWR.n107 VAPWR.n80 184.847
R617 VAPWR.n82 VAPWR.n80 184.847
R618 VAPWR.n59 VAPWR.n5 172.655
R619 VAPWR.n111 VAPWR.n74 172.655
R620 VAPWR.n55 VAPWR.t12 167.41
R621 VAPWR.n79 VAPWR.t15 167.41
R622 VAPWR.n120 VAPWR.t8 167.251
R623 VAPWR.n68 VAPWR.t16 167.141
R624 VAPWR.n60 VAPWR.n59 160.495
R625 VAPWR.n112 VAPWR.n111 160.495
R626 VAPWR.n107 VAPWR.n81 146.25
R627 VAPWR.n83 VAPWR.n82 146.25
R628 VAPWR.n106 VAPWR.n87 97.5005
R629 VAPWR.n84 VAPWR.n80 97.5005
R630 VAPWR.n105 VAPWR.t4 82.8472
R631 VAPWR.t9 VAPWR.t11 81.0585
R632 VAPWR.t13 VAPWR.t7 81.0585
R633 VAPWR.n85 VAPWR.n83 72.5386
R634 VAPWR.n86 VAPWR.n81 72.5386
R635 VAPWR.n86 VAPWR.t3 66.988
R636 VAPWR.t3 VAPWR.n85 66.988
R637 VAPWR.n63 VAPWR.n61 34.0449
R638 VAPWR.n115 VAPWR.n113 34.0449
R639 VAPWR.n62 VAPWR.n3 23.1255
R640 VAPWR.n63 VAPWR.n62 23.1255
R641 VAPWR.n65 VAPWR.n64 23.1255
R642 VAPWR.n114 VAPWR.n72 23.1255
R643 VAPWR.n115 VAPWR.n114 23.1255
R644 VAPWR.n117 VAPWR.n116 23.1255
R645 VAPWR.t9 VAPWR.n61 21.1116
R646 VAPWR.t13 VAPWR.n113 21.1116
R647 VAPWR.n43 VAPWR.n37 14.2313
R648 VAPWR.n44 VAPWR.n43 14.2313
R649 VAPWR.n48 VAPWR.n47 14.2313
R650 VAPWR.n47 VAPWR.n46 14.2313
R651 VAPWR.n26 VAPWR.n20 14.2313
R652 VAPWR.n27 VAPWR.n26 14.2313
R653 VAPWR.n31 VAPWR.n30 14.2313
R654 VAPWR.n30 VAPWR.n29 14.2313
R655 VAPWR.n15 VAPWR.n14 14.2313
R656 VAPWR.n14 VAPWR.n13 14.2313
R657 VAPWR.n58 VAPWR.n57 14.2313
R658 VAPWR.n59 VAPWR.n58 14.2313
R659 VAPWR.n95 VAPWR.n94 14.2313
R660 VAPWR.n94 VAPWR.n93 14.2313
R661 VAPWR.n110 VAPWR.n109 14.2313
R662 VAPWR.n111 VAPWR.n110 14.2313
R663 VAPWR.n41 VAPWR.n40 12.3338
R664 VAPWR.n42 VAPWR.n41 12.3338
R665 VAPWR.n49 VAPWR.n38 12.3338
R666 VAPWR.n45 VAPWR.n38 12.3338
R667 VAPWR.n24 VAPWR.n23 12.3338
R668 VAPWR.n25 VAPWR.n24 12.3338
R669 VAPWR.n32 VAPWR.n21 12.3338
R670 VAPWR.n28 VAPWR.n21 12.3338
R671 VAPWR.n8 VAPWR.n6 12.3338
R672 VAPWR.n11 VAPWR.n6 12.3338
R673 VAPWR.n9 VAPWR.n7 12.3338
R674 VAPWR.n12 VAPWR.n7 12.3338
R675 VAPWR.n78 VAPWR.n76 12.3338
R676 VAPWR.n92 VAPWR.n76 12.3338
R677 VAPWR.n77 VAPWR.n75 12.3338
R678 VAPWR.n91 VAPWR.n75 12.3338
R679 VAPWR.n66 VAPWR.n4 7.70883
R680 VAPWR.n60 VAPWR.n4 7.70883
R681 VAPWR.n118 VAPWR.n73 7.70883
R682 VAPWR.n112 VAPWR.n73 7.70883
R683 VAPWR.n125 VAPWR 4.11654
R684 VAPWR.n126 VAPWR 4.06671
R685 VAPWR.n123 VAPWR 3.16715
R686 VAPWR.n123 VAPWR 3.13288
R687 VAPWR.n39 VAPWR.n35 2.77496
R688 VAPWR.n39 VAPWR.n36 2.77496
R689 VAPWR.n50 VAPWR.n36 2.77496
R690 VAPWR.n22 VAPWR.n18 2.77496
R691 VAPWR.n22 VAPWR.n19 2.77496
R692 VAPWR.n33 VAPWR.n19 2.77496
R693 VAPWR.n16 VAPWR.n10 2.77496
R694 VAPWR.n17 VAPWR.n16 2.77496
R695 VAPWR.n98 VAPWR.n82 2.3255
R696 VAPWR.n108 VAPWR.n107 2.3255
R697 VAPWR.n54 VAPWR.n3 2.1216
R698 VAPWR.n89 VAPWR.n72 2.09672
R699 VAPWR.n52 VAPWR.n34 1.88425
R700 VAPWR.n106 VAPWR.n105 1.5505
R701 VAPWR.n10 VAPWR 1.40267
R702 VAPWR.n53 VAPWR.n52 1.37675
R703 VAPWR.n96 VAPWR.n95 1.32345
R704 VAPWR.n53 VAPWR.n17 1.23691
R705 VAPWR.n51 VAPWR.n50 1.22254
R706 VAPWR.n34 VAPWR.n33 1.22254
R707 VAPWR.n65 VAPWR.n1 1.163
R708 VAPWR.n117 VAPWR.n71 1.163
R709 VAPWR.n124 VAPWR.n123 1.07737
R710 VAPWR.n51 VAPWR.n35 0.894522
R711 VAPWR.n34 VAPWR.n18 0.894522
R712 VAPWR.n48 VAPWR.n35 0.845955
R713 VAPWR.n37 VAPWR.n36 0.845955
R714 VAPWR.n31 VAPWR.n18 0.845955
R715 VAPWR.n20 VAPWR.n19 0.845955
R716 VAPWR.n16 VAPWR.n15 0.845955
R717 VAPWR.n57 VAPWR.n56 0.845955
R718 VAPWR.n109 VAPWR.n108 0.845955
R719 VAPWR.t11 VAPWR.n63 0.81108
R720 VAPWR.t7 VAPWR.n115 0.81108
R721 VAPWR.n104 VAPWR.n103 0.797375
R722 VAPWR.n40 VAPWR.n39 0.664786
R723 VAPWR.n50 VAPWR.n49 0.664786
R724 VAPWR.n23 VAPWR.n22 0.664786
R725 VAPWR.n33 VAPWR.n32 0.664786
R726 VAPWR.n10 VAPWR.n9 0.664786
R727 VAPWR.n17 VAPWR.n8 0.664786
R728 VAPWR.n101 VAPWR.n78 0.664786
R729 VAPWR.n90 VAPWR.n77 0.664786
R730 VAPWR.n52 VAPWR.n51 0.5005
R731 VAPWR VAPWR.n126 0.491143
R732 VAPWR VAPWR.n88 0.490083
R733 VAPWR.n70 VAPWR.n1 0.448327
R734 VAPWR.n67 VAPWR.n66 0.404848
R735 VAPWR.n119 VAPWR.n118 0.404848
R736 VAPWR.n98 VAPWR.n97 0.3455
R737 VAPWR.n68 VAPWR.n0 0.313
R738 VAPWR.n125 VAPWR.n124 0.2968
R739 VAPWR.n103 VAPWR.n102 0.203625
R740 VAPWR.n96 VAPWR.n90 0.198256
R741 VAPWR.n70 VAPWR.n0 0.188
R742 VAPWR.n55 VAPWR.n54 0.179291
R743 VAPWR.n99 VAPWR.n98 0.163
R744 VAPWR.n56 VAPWR.n2 0.157262
R745 VAPWR.n119 VAPWR 0.152375
R746 VAPWR.n69 VAPWR.n68 0.143
R747 VAPWR.n101 VAPWR.n100 0.14175
R748 VAPWR.n70 VAPWR.n69 0.140949
R749 VAPWR VAPWR.n2 0.136533
R750 VAPWR.n104 VAPWR.n88 0.130708
R751 VAPWR VAPWR.n121 0.123855
R752 VAPWR VAPWR.n70 0.105837
R753 VAPWR.n90 VAPWR.n89 0.0951602
R754 VAPWR.n103 VAPWR.n101 0.0905
R755 VAPWR.n89 VAPWR.n79 0.0695895
R756 VAPWR.n121 VAPWR.n120 0.0690307
R757 VAPWR.n124 VAPWR 0.0651875
R758 VAPWR.n67 VAPWR.n2 0.062375
R759 VAPWR.n105 VAPWR 0.0568725
R760 VAPWR.n100 VAPWR.n99 0.0544216
R761 VAPWR.n122 VAPWR.n71 0.0533274
R762 VAPWR.n97 VAPWR 0.043
R763 VAPWR.n100 VAPWR 0.0364477
R764 VAPWR.n105 VAPWR 0.0364477
R765 VAPWR.n120 VAPWR.n119 0.033625
R766 VAPWR.n99 VAPWR.n96 0.0305
R767 VAPWR.n102 VAPWR 0.029875
R768 VAPWR.n56 VAPWR.n55 0.0297008
R769 VAPWR VAPWR.n122 0.0235263
R770 VAPWR VAPWR.n88 0.0212668
R771 VAPWR.n88 VAPWR 0.01927
R772 VAPWR VAPWR.n104 0.0184739
R773 VAPWR.n102 VAPWR 0.0152764
R774 VAPWR.n108 VAPWR.n79 0.0118818
R775 VAPWR.n108 VAPWR 0.00728914
R776 VAPWR.n122 VAPWR 0.00488596
R777 VAPWR.n54 VAPWR.n53 0.00425
R778 VAPWR.n126 VAPWR.n125 0.0033356
R779 VAPWR.n69 VAPWR.n67 0.002375
R780 flash_0.x2.clkb flash_0.x2.clkb.t0 167.038
R781 flash_0.x2.clkb flash_0.x2.clkb.t1 87.4292
R782 clk.n1 clk.t2 54.3383
R783 clk.n0 clk.t0 54.3383
R784 clk.n1 clk.t3 53.1307
R785 clk.n0 clk.t1 53.1307
R786 clk.n3 clk 39.2423
R787 clk.n3 clk.n2 9.04175
R788 clk.n2 clk 7.02925
R789 clk.n2 clk 3.72425
R790 clk clk.n1 0.2455
R791 clk clk.n0 0.2455
R792 clk clk.n3 0.078
R793 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t1 649.691
R794 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t2 227.442
R795 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t0 227.361
R796 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t5 216.731
R797 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t6 216.731
R798 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t3 216.731
R799 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t4 216.731
R800 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t7 216.731
R801 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t8 216.731
R802 ui_in[1].n0 ui_in[1].t17 207.43
R803 ui_in[1].n1 ui_in[1].t10 207.43
R804 ui_in[1].n2 ui_in[1].t12 207.43
R805 ui_in[1].n3 ui_in[1].t13 207.43
R806 ui_in[1].n4 ui_in[1].t15 207.43
R807 ui_in[1].n5 ui_in[1].t2 207.43
R808 ui_in[1].n26 ui_in[1].n23 123.867
R809 ui_in[1].n25 ui_in[1] 50.8126
R810 ui_in[1].n15 ui_in[1] 50.8126
R811 ui_in[1] ui_in[1].n1 48.5522
R812 ui_in[1] ui_in[1].n3 48.5522
R813 ui_in[1].n6 ui_in[1].n5 47.7953
R814 ui_in[1].n6 ui_in[1].n2 32.1435
R815 ui_in[1].n8 ui_in[1] 29.9794
R816 ui_in[1].n10 ui_in[1] 29.9794
R817 ui_in[1].n21 ui_in[1] 29.418
R818 ui_in[1].n18 ui_in[1] 29.418
R819 ui_in[1].n27 ui_in[1] 22.2876
R820 ui_in[1].n25 ui_in[1].n24 19.0005
R821 ui_in[1].n21 ui_in[1].n20 19.0005
R822 ui_in[1].n18 ui_in[1].n17 19.0005
R823 ui_in[1].n15 ui_in[1].n14 19.0005
R824 ui_in[1].n8 ui_in[1].n7 19.0005
R825 ui_in[1].n10 ui_in[1].n9 19.0005
R826 ui_in[1] ui_in[1].n0 13.6833
R827 ui_in[1] ui_in[1].n4 13.6833
R828 ui_in[1].n20 ui_in[1].t9 12.0505
R829 ui_in[1].n20 ui_in[1].t6 12.0505
R830 ui_in[1].n17 ui_in[1].t11 12.0505
R831 ui_in[1].n17 ui_in[1].t8 12.0505
R832 ui_in[1].n7 ui_in[1].t5 12.0505
R833 ui_in[1].n7 ui_in[1].t0 12.0505
R834 ui_in[1].n9 ui_in[1].t16 12.0505
R835 ui_in[1].n9 ui_in[1].t14 12.0505
R836 ui_in[1].n27 ui_in[1] 8.72144
R837 ui_in[1].n24 ui_in[1].t3 8.4355
R838 ui_in[1].n24 ui_in[1].t1 8.4355
R839 ui_in[1].n14 ui_in[1].t7 8.4355
R840 ui_in[1].n14 ui_in[1].t4 8.4355
R841 ui_in[1] ui_in[1].n26 4.94473
R842 ui_in[1].n13 ui_in[1].n12 4.5005
R843 ui_in[1].n2 ui_in[1] 3.75222
R844 ui_in[1].n1 ui_in[1] 3.75222
R845 ui_in[1].n0 ui_in[1] 3.75222
R846 ui_in[1].n5 ui_in[1] 3.75222
R847 ui_in[1].n4 ui_in[1] 3.75222
R848 ui_in[1].n3 ui_in[1] 3.75222
R849 ui_in[1].n28 ui_in[1].n13 3.61982
R850 ui_in[1].n11 ui_in[1].n8 2.96269
R851 ui_in[1].n12 ui_in[1].n6 1.69929
R852 ui_in[1].n16 ui_in[1].n15 1.59032
R853 ui_in[1].n22 ui_in[1].n19 1.42722
R854 ui_in[1].n19 ui_in[1].n18 1.32907
R855 ui_in[1].n22 ui_in[1].n21 1.32907
R856 ui_in[1].n26 ui_in[1].n25 1.32907
R857 ui_in[1].n11 ui_in[1].n10 1.32907
R858 ui_in[1].n23 ui_in[1].n16 1.29347
R859 ui_in[1].n12 ui_in[1].n11 0.48697
R860 ui_in[1].n19 ui_in[1].n16 0.25925
R861 ui_in[1].n23 ui_in[1].n22 0.25925
R862 ui_in[1].n13 ui_in[1] 0.0611061
R863 ui_in[1].n28 ui_in[1].n27 0.039875
R864 ui_in[1] ui_in[1].n28 0.0214375
R865 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t3 669.481
R866 flash_0.x4.neg_en_b.n0 flash_0.x4.neg_en_b.t0 669.481
R867 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t1 218.06
R868 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t2 218.06
R869 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t4 211.017
R870 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t6 208.394
R871 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t9 208.394
R872 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t5 207.43
R873 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t7 207.43
R874 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t8 207.43
R875 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.n0 50.3013
R876 flash_0.x4.neg_en_b.n0 flash_0.x4.neg_en_b 29.0914
R877 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t5 649.773
R878 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t1 649.691
R879 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.n1 594.383
R880 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.n2 594.301
R881 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t0 227.361
R882 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t8 216.731
R883 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t14 216.731
R884 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t13 216.731
R885 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t9 105.956
R886 flash_0.x4.neg_mid_b.n0 flash_0.x4.neg_mid_b 103.529
R887 flash_0.x4.neg_mid_b.t8 flash_0.x4.neg_mid_b.t7 101.221
R888 flash_0.x4.neg_mid_b.t14 flash_0.x4.neg_mid_b.t12 101.221
R889 flash_0.x4.neg_mid_b.t13 flash_0.x4.neg_mid_b.t11 101.221
R890 flash_0.x4.neg_mid_b.n2 flash_0.x4.neg_mid_b.t2 55.3905
R891 flash_0.x4.neg_mid_b.n2 flash_0.x4.neg_mid_b.t6 55.3905
R892 flash_0.x4.neg_mid_b.n1 flash_0.x4.neg_mid_b.t3 55.3905
R893 flash_0.x4.neg_mid_b.n1 flash_0.x4.neg_mid_b.t4 55.3905
R894 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.n0 23.6062
R895 flash_0.x4.neg_mid_b.n0 flash_0.x4.neg_mid_b.t10 22.3887
R896 flash_0.x4.VOUT flash_0.x4.VOUT.t3 649.691
R897 flash_0.x4.VOUT flash_0.x4.VOUT.t10 649.691
R898 flash_0.x4.VOUT flash_0.x4.VOUT.t8 649.691
R899 flash_0.x4.VOUT flash_0.x4.VOUT.t1 649.691
R900 flash_0.x4.VOUT flash_0.x4.VOUT.n0 594.383
R901 flash_0.x4.VOUT flash_0.x4.VOUT.n2 594.301
R902 flash_0.x4.VOUT flash_0.x4.VOUT.n3 594.301
R903 flash_0.x4.VOUT flash_0.x4.VOUT.n1 594.301
R904 flash_0.x4.VOUT flash_0.x4.VOUT.t4 227.431
R905 flash_0.x4.VOUT flash_0.x4.VOUT.t0 227.361
R906 flash_0.x4.VOUT flash_0.x4.VOUT.t14 149.423
R907 flash_0.x4.VOUT.n2 flash_0.x4.VOUT.t2 55.3905
R908 flash_0.x4.VOUT.n2 flash_0.x4.VOUT.t12 55.3905
R909 flash_0.x4.VOUT.n3 flash_0.x4.VOUT.t13 55.3905
R910 flash_0.x4.VOUT.n3 flash_0.x4.VOUT.t5 55.3905
R911 flash_0.x4.VOUT.n1 flash_0.x4.VOUT.t11 55.3905
R912 flash_0.x4.VOUT.n1 flash_0.x4.VOUT.t9 55.3905
R913 flash_0.x4.VOUT.n0 flash_0.x4.VOUT.t7 55.3905
R914 flash_0.x4.VOUT.n0 flash_0.x4.VOUT.t6 55.3905
R915 flash_0.x4.dcgint.n0 flash_0.x4.dcgint.t8 644.461
R916 flash_0.x4.dcgint.n5 flash_0.x4.dcgint.t6 640.39
R917 flash_0.x4.dcgint.n3 flash_0.x4.dcgint.n1 605.365
R918 flash_0.x4.dcgint.n3 flash_0.x4.dcgint.n2 605.365
R919 flash_0.x4.dcgint.n4 flash_0.x4.dcgint.t5 477.228
R920 flash_0.x4.dcgint.t5 flash_0.x4.dcgint.t3 339.594
R921 flash_0.x4.dcgint.t3 flash_0.x4.dcgint.t9 339.594
R922 flash_0.x4.dcgint flash_0.x4.dcgint.t2 227.361
R923 flash_0.x4.dcgint flash_0.x4.dcgint.t1 227.361
R924 flash_0.x4.dcgint flash_0.x4.dcgint.t0 227.361
R925 flash_0.x4.dcgint.n4 flash_0.x4.dcgint.n3 69.5657
R926 flash_0.x4.dcgint.n1 flash_0.x4.dcgint.t4 55.3905
R927 flash_0.x4.dcgint.n1 flash_0.x4.dcgint.t10 55.3905
R928 flash_0.x4.dcgint.n2 flash_0.x4.dcgint.t7 55.3905
R929 flash_0.x4.dcgint.n2 flash_0.x4.dcgint.t11 55.3905
R930 flash_0.x4.dcgint.n6 flash_0.x4.dcgint.n5 9.3005
R931 flash_0.x4.dcgint.n5 flash_0.x4.dcgint.n4 8.9605
R932 flash_0.x4.dcgint flash_0.x4.dcgint.n6 7.52362
R933 flash_0.x4.dcgint.n6 flash_0.x4.dcgint.n0 1.14684
R934 flash_0.x4.dcgint.n4 flash_0.x4.dcgint.n0 1.0086
R935 flash_0.x7.pos_en_b.n1 flash_0.x7.pos_en_b.t1 669.481
R936 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b.t0 669.481
R937 flash_0.x7.pos_en_b flash_0.x7.pos_en_b.t2 218.06
R938 flash_0.x7.pos_en_b flash_0.x7.pos_en_b.t3 218.06
R939 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b.t6 65.4032
R940 flash_0.x7.pos_en_b.t6 flash_0.x7.pos_en_b 56.2429
R941 flash_0.x7.pos_en_b.t6 flash_0.x7.pos_en_b 56.2429
R942 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b 50.8126
R943 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b 50.8126
R944 flash_0.x7.pos_en_b flash_0.x7.pos_en_b.n1 29.0914
R945 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b 29.0914
R946 flash_0.x7.pos_en_b.n1 flash_0.x7.pos_en_b.n0 28.2591
R947 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b.t4 27.4355
R948 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b.t5 27.4355
R949 VDPWR.n103 VDPWR.n89 5586
R950 VDPWR.n103 VDPWR.n90 5586
R951 VDPWR.n98 VDPWR.n90 5586
R952 VDPWR.n98 VDPWR.n89 5586
R953 VDPWR.n148 VDPWR.n134 5586
R954 VDPWR.n148 VDPWR.n135 5586
R955 VDPWR.n143 VDPWR.n135 5586
R956 VDPWR.n143 VDPWR.n134 5586
R957 VDPWR.n49 VDPWR.n48 4689.72
R958 VDPWR.n46 VDPWR.n44 4689.72
R959 VDPWR.n99 VDPWR.n91 4509.29
R960 VDPWR.n144 VDPWR.n136 4509.29
R961 VDPWR.n102 VDPWR.n91 4506
R962 VDPWR.n147 VDPWR.n136 4506
R963 VDPWR.n63 VDPWR.n56 2442.35
R964 VDPWR.n60 VDPWR.n57 2442.35
R965 VDPWR.n80 VDPWR.n73 2442.35
R966 VDPWR.n77 VDPWR.n74 2442.35
R967 VDPWR.n102 VDPWR.t6 2271.78
R968 VDPWR.n147 VDPWR.t31 2271.78
R969 VDPWR.n49 VDPWR.n43 1828.1
R970 VDPWR.n47 VDPWR.n46 1828.1
R971 VDPWR.t10 VDPWR.t37 1429.17
R972 VDPWR.t35 VDPWR.t0 1429.17
R973 VDPWR.t6 VDPWR.n101 1226.56
R974 VDPWR.t31 VDPWR.n146 1226.56
R975 VDPWR.n45 VDPWR.n41 902.777
R976 VDPWR.n45 VDPWR.n42 902.777
R977 VDPWR.n50 VDPWR.n42 881.453
R978 VDPWR.n51 VDPWR.n41 879.466
R979 VDPWR.n52 VDPWR.t54 649.831
R980 VDPWR.n104 VDPWR.n88 627.201
R981 VDPWR.n97 VDPWR.n87 627.201
R982 VDPWR.n149 VDPWR.n133 627.201
R983 VDPWR.n142 VDPWR.n132 627.201
R984 VDPWR.n123 VDPWR.n122 585
R985 VDPWR.n118 VDPWR.n117 585
R986 VDPWR.n113 VDPWR.n112 585
R987 VDPWR.n121 VDPWR.n120 585
R988 VDPWR.n116 VDPWR.n115 585
R989 VDPWR.n111 VDPWR.n110 585
R990 VDPWR.n22 VDPWR.n21 585
R991 VDPWR.n17 VDPWR.n16 585
R992 VDPWR.n12 VDPWR.n11 585
R993 VDPWR.n20 VDPWR.n19 585
R994 VDPWR.n15 VDPWR.n14 585
R995 VDPWR.n10 VDPWR.n9 585
R996 VDPWR.n61 VDPWR.n56 535.419
R997 VDPWR.n62 VDPWR.n57 535.419
R998 VDPWR.n78 VDPWR.n73 535.419
R999 VDPWR.n79 VDPWR.n74 535.419
R1000 VDPWR.n105 VDPWR.n104 525.553
R1001 VDPWR.n150 VDPWR.n149 525.553
R1002 VDPWR.n96 VDPWR.n88 492.048
R1003 VDPWR.n141 VDPWR.n133 492.048
R1004 VDPWR.n101 VDPWR.t10 394.779
R1005 VDPWR.n146 VDPWR.t35 394.779
R1006 VDPWR.n107 VDPWR.n85 297.151
R1007 VDPWR.n127 VDPWR.n126 297.151
R1008 VDPWR.n26 VDPWR.n25 297.151
R1009 VDPWR.n152 VDPWR.n130 297.151
R1010 VDPWR.n100 VDPWR.t27 272.363
R1011 VDPWR.n145 VDPWR.t42 272.363
R1012 VDPWR.n59 VDPWR.n55 260.519
R1013 VDPWR.n64 VDPWR.n55 260.519
R1014 VDPWR.n76 VDPWR.n72 260.519
R1015 VDPWR.n81 VDPWR.n72 260.519
R1016 VDPWR.n59 VDPWR.n58 232.66
R1017 VDPWR.n65 VDPWR.n64 232.66
R1018 VDPWR.n76 VDPWR.n75 232.66
R1019 VDPWR.n82 VDPWR.n81 232.66
R1020 VDPWR.n53 VDPWR.t13 228.215
R1021 VDPWR.n70 VDPWR.t45 228.215
R1022 VDPWR VDPWR.t69 216.822
R1023 VDPWR VDPWR.t62 216.822
R1024 VDPWR.n35 VDPWR.t58 216.731
R1025 VDPWR.n32 VDPWR.t63 216.731
R1026 VDPWR.n33 VDPWR.t64 216.731
R1027 VDPWR.n30 VDPWR.t60 216.731
R1028 VDPWR.n29 VDPWR.t67 216.731
R1029 VDPWR.n6 VDPWR.t65 216.731
R1030 VDPWR.n3 VDPWR.t70 216.731
R1031 VDPWR.n4 VDPWR.t71 216.731
R1032 VDPWR.n1 VDPWR.t72 216.731
R1033 VDPWR.n0 VDPWR.t73 216.731
R1034 VDPWR.t39 VDPWR.t29 172.133
R1035 VDPWR.t33 VDPWR.t25 172.133
R1036 VDPWR.t21 VDPWR.t33 172.133
R1037 VDPWR.t27 VDPWR.t21 172.133
R1038 VDPWR.t2 VDPWR.t14 172.133
R1039 VDPWR.t16 VDPWR.t4 172.133
R1040 VDPWR.t8 VDPWR.t16 172.133
R1041 VDPWR.t42 VDPWR.t8 172.133
R1042 VDPWR.n85 VDPWR.t11 160.44
R1043 VDPWR.n85 VDPWR.t7 160.44
R1044 VDPWR.n126 VDPWR.t24 160.44
R1045 VDPWR.n126 VDPWR.t38 160.44
R1046 VDPWR.n25 VDPWR.t20 160.44
R1047 VDPWR.n25 VDPWR.t1 160.44
R1048 VDPWR.n130 VDPWR.t36 160.44
R1049 VDPWR.n130 VDPWR.t32 160.44
R1050 VDPWR.n97 VDPWR.n96 135.154
R1051 VDPWR.n142 VDPWR.n141 135.154
R1052 VDPWR.t23 VDPWR.t39 135.093
R1053 VDPWR.t19 VDPWR.t2 135.093
R1054 VDPWR.n93 VDPWR 106.918
R1055 VDPWR.n138 VDPWR 106.918
R1056 VDPWR.n105 VDPWR.n87 101.647
R1057 VDPWR.n150 VDPWR.n132 101.647
R1058 VDPWR.n100 VDPWR.n99 57.7708
R1059 VDPWR.n145 VDPWR.n144 57.7708
R1060 VDPWR.n122 VDPWR.t22 55.3905
R1061 VDPWR.n122 VDPWR.t50 55.3905
R1062 VDPWR.n117 VDPWR.t48 55.3905
R1063 VDPWR.n117 VDPWR.t34 55.3905
R1064 VDPWR.n112 VDPWR.t30 55.3905
R1065 VDPWR.n112 VDPWR.t47 55.3905
R1066 VDPWR.n120 VDPWR.t49 55.3905
R1067 VDPWR.n120 VDPWR.t28 55.3905
R1068 VDPWR.n115 VDPWR.t26 55.3905
R1069 VDPWR.n115 VDPWR.t46 55.3905
R1070 VDPWR.n110 VDPWR.t51 55.3905
R1071 VDPWR.n110 VDPWR.t40 55.3905
R1072 VDPWR.n21 VDPWR.t9 55.3905
R1073 VDPWR.n21 VDPWR.t56 55.3905
R1074 VDPWR.n16 VDPWR.t5 55.3905
R1075 VDPWR.n16 VDPWR.t17 55.3905
R1076 VDPWR.n11 VDPWR.t57 55.3905
R1077 VDPWR.n11 VDPWR.t52 55.3905
R1078 VDPWR.n19 VDPWR.t55 55.3905
R1079 VDPWR.n19 VDPWR.t43 55.3905
R1080 VDPWR.n14 VDPWR.t18 55.3905
R1081 VDPWR.n14 VDPWR.t41 55.3905
R1082 VDPWR.n9 VDPWR.t15 55.3905
R1083 VDPWR.n9 VDPWR.t3 55.3905
R1084 VDPWR.t25 VDPWR.t23 37.0418
R1085 VDPWR.t4 VDPWR.t19 37.0418
R1086 VDPWR.n46 VDPWR.n45 37.0005
R1087 VDPWR.n50 VDPWR.n49 37.0005
R1088 VDPWR.n57 VDPWR.n55 30.8338
R1089 VDPWR.n56 VDPWR.n54 30.8338
R1090 VDPWR.n74 VDPWR.n72 30.8338
R1091 VDPWR.n73 VDPWR.n71 30.8338
R1092 VDPWR.n58 VDPWR.n54 27.8593
R1093 VDPWR.n65 VDPWR.n54 27.8593
R1094 VDPWR.n75 VDPWR.n71 27.8593
R1095 VDPWR.n82 VDPWR.n71 27.8593
R1096 VDPWR.n93 VDPWR.n92 19.0005
R1097 VDPWR.n138 VDPWR.n137 19.0005
R1098 VDPWR.n60 VDPWR.n59 16.8187
R1099 VDPWR.n64 VDPWR.n63 16.8187
R1100 VDPWR.n77 VDPWR.n76 16.8187
R1101 VDPWR.n81 VDPWR.n80 16.8187
R1102 VDPWR.n123 VDPWR 14.3064
R1103 VDPWR.n118 VDPWR 14.3064
R1104 VDPWR.n113 VDPWR 14.3064
R1105 VDPWR.n121 VDPWR 14.3064
R1106 VDPWR.n116 VDPWR 14.3064
R1107 VDPWR.n111 VDPWR 14.3064
R1108 VDPWR.n22 VDPWR 14.3064
R1109 VDPWR.n17 VDPWR 14.3064
R1110 VDPWR.n12 VDPWR 14.3064
R1111 VDPWR.n20 VDPWR 14.3064
R1112 VDPWR.n15 VDPWR 14.3064
R1113 VDPWR.n10 VDPWR 14.3064
R1114 VDPWR.n124 VDPWR.n123 13.8019
R1115 VDPWR.n119 VDPWR.n118 13.8019
R1116 VDPWR.n114 VDPWR.n113 13.8019
R1117 VDPWR.n124 VDPWR.n121 13.8019
R1118 VDPWR.n119 VDPWR.n116 13.8019
R1119 VDPWR.n114 VDPWR.n111 13.8019
R1120 VDPWR.n23 VDPWR.n22 13.8019
R1121 VDPWR.n18 VDPWR.n17 13.8019
R1122 VDPWR.n13 VDPWR.n12 13.8019
R1123 VDPWR.n23 VDPWR.n20 13.8019
R1124 VDPWR.n18 VDPWR.n15 13.8019
R1125 VDPWR.n13 VDPWR.n10 13.8019
R1126 VDPWR.n61 VDPWR.n60 13.0425
R1127 VDPWR.n63 VDPWR.n62 13.0425
R1128 VDPWR.n78 VDPWR.n77 13.0425
R1129 VDPWR.n80 VDPWR.n79 13.0425
R1130 VDPWR.t37 VDPWR.n100 10.895
R1131 VDPWR.t0 VDPWR.n145 10.895
R1132 VDPWR.n104 VDPWR.n103 10.2783
R1133 VDPWR.n103 VDPWR.n102 10.2783
R1134 VDPWR.n98 VDPWR.n97 10.2783
R1135 VDPWR.n99 VDPWR.n98 10.2783
R1136 VDPWR.n149 VDPWR.n148 10.2783
R1137 VDPWR.n148 VDPWR.n147 10.2783
R1138 VDPWR.n143 VDPWR.n142 10.2783
R1139 VDPWR.n144 VDPWR.n143 10.2783
R1140 VDPWR.n84 VDPWR.n83 9.74376
R1141 VDPWR.n58 VDPWR.n53 9.35589
R1142 VDPWR.n75 VDPWR.n70 9.35589
R1143 VDPWR VDPWR.n65 9.33194
R1144 VDPWR VDPWR.n82 9.33194
R1145 VDPWR.n92 VDPWR.t61 8.4355
R1146 VDPWR.n92 VDPWR.t59 8.4355
R1147 VDPWR.n137 VDPWR.t68 8.4355
R1148 VDPWR.n137 VDPWR.t66 8.4355
R1149 VDPWR.n89 VDPWR.n88 6.37981
R1150 VDPWR.n91 VDPWR.n89 6.37981
R1151 VDPWR.n90 VDPWR.n87 6.37981
R1152 VDPWR.n101 VDPWR.n90 6.37981
R1153 VDPWR.n134 VDPWR.n133 6.37981
R1154 VDPWR.n136 VDPWR.n134 6.37981
R1155 VDPWR.n135 VDPWR.n132 6.37981
R1156 VDPWR.n146 VDPWR.n135 6.37981
R1157 VDPWR.n67 VDPWR.n52 5.59737
R1158 VDPWR.n94 VDPWR.n86 4.51137
R1159 VDPWR.n139 VDPWR.n131 4.51137
R1160 VDPWR.n153 VDPWR.n152 3.96097
R1161 VDPWR.n108 VDPWR.n107 3.9605
R1162 VDPWR.n96 VDPWR.n95 3.88885
R1163 VDPWR.n141 VDPWR.n140 3.88885
R1164 VDPWR.n39 VDPWR 3.84311
R1165 VDPWR.n109 VDPWR.n38 3.79423
R1166 VDPWR.n106 VDPWR.n86 3.7551
R1167 VDPWR.n151 VDPWR.n131 3.7551
R1168 VDPWR.n62 VDPWR.t12 3.68792
R1169 VDPWR.t12 VDPWR.n61 3.68792
R1170 VDPWR.n79 VDPWR.t44 3.68792
R1171 VDPWR.t44 VDPWR.n78 3.68792
R1172 VDPWR.n44 VDPWR.n41 3.03329
R1173 VDPWR.n48 VDPWR.n42 3.03329
R1174 VDPWR.n95 VDPWR.n93 2.3749
R1175 VDPWR.n140 VDPWR.n138 2.3749
R1176 VDPWR.n27 VDPWR.n26 2.25658
R1177 VDPWR.n128 VDPWR.n127 2.2555
R1178 VDPWR.n37 VDPWR.n36 2.2505
R1179 VDPWR.n8 VDPWR.n7 2.2505
R1180 VDPWR.n155 VDPWR.n154 2.08954
R1181 VDPWR.n154 VDPWR.n27 1.8913
R1182 VDPWR.n52 VDPWR.n51 1.8605
R1183 VDPWR.n44 VDPWR.n43 1.85038
R1184 VDPWR.n48 VDPWR.n47 1.85038
R1185 VDPWR.n129 VDPWR.n128 1.7055
R1186 VDPWR.n68 VDPWR.n67 1.43592
R1187 VDPWR.n84 VDPWR.n69 1.29333
R1188 VDPWR.n47 VDPWR.t53 1.18321
R1189 VDPWR.t53 VDPWR.n43 1.18321
R1190 VDPWR.n51 VDPWR.n50 1.0245
R1191 VDPWR.n95 VDPWR.n94 0.813
R1192 VDPWR.n140 VDPWR.n139 0.813
R1193 VDPWR.n108 VDPWR.n84 0.683034
R1194 VDPWR.n156 VDPWR 0.59425
R1195 VDPWR.n104 VDPWR.n86 0.547559
R1196 VDPWR.n149 VDPWR.n131 0.547559
R1197 VDPWR.n67 VDPWR.n66 0.53175
R1198 VDPWR.n69 VDPWR.n68 0.486785
R1199 VDPWR.n153 VDPWR.n129 0.475641
R1200 VDPWR.n106 VDPWR.n105 0.4655
R1201 VDPWR.n151 VDPWR.n150 0.4655
R1202 VDPWR.n94 VDPWR.n88 0.344944
R1203 VDPWR.n139 VDPWR.n133 0.344944
R1204 VDPWR.n28 VDPWR 0.339786
R1205 VDPWR VDPWR.n33 0.337457
R1206 VDPWR VDPWR.n32 0.337457
R1207 VDPWR.n29 VDPWR 0.337457
R1208 VDPWR.n30 VDPWR 0.337457
R1209 VDPWR VDPWR.n4 0.337457
R1210 VDPWR VDPWR.n3 0.337457
R1211 VDPWR.n0 VDPWR 0.337457
R1212 VDPWR.n1 VDPWR 0.337457
R1213 VDPWR.n38 VDPWR 0.326693
R1214 VDPWR.n8 VDPWR 0.317148
R1215 VDPWR.n27 VDPWR.n24 0.201021
R1216 VDPWR.n129 VDPWR.n109 0.186297
R1217 VDPWR.n128 VDPWR.n125 0.182167
R1218 VDPWR.n40 VDPWR.n39 0.171
R1219 VDPWR.n36 VDPWR.n35 0.122211
R1220 VDPWR.n7 VDPWR.n6 0.122211
R1221 VDPWR.n127 VDPWR 0.102773
R1222 VDPWR.n26 VDPWR 0.102773
R1223 VDPWR.n154 VDPWR.n153 0.0952344
R1224 VDPWR.n37 VDPWR.n28 0.0935233
R1225 VDPWR.n33 VDPWR 0.0928913
R1226 VDPWR.n32 VDPWR 0.0928913
R1227 VDPWR VDPWR.n29 0.0928913
R1228 VDPWR.n4 VDPWR 0.0928913
R1229 VDPWR.n3 VDPWR 0.0928913
R1230 VDPWR VDPWR.n0 0.0928913
R1231 VDPWR.n156 VDPWR.n155 0.0928913
R1232 VDPWR.n109 VDPWR.n108 0.0928088
R1233 VDPWR.n119 VDPWR.n114 0.0902727
R1234 VDPWR.n18 VDPWR.n13 0.0902727
R1235 VDPWR.n36 VDPWR 0.0827368
R1236 VDPWR.n7 VDPWR 0.0827368
R1237 VDPWR.n34 VDPWR 0.0820217
R1238 VDPWR.n5 VDPWR 0.0820217
R1239 VDPWR.n125 VDPWR.n119 0.0772045
R1240 VDPWR.n24 VDPWR.n18 0.0772045
R1241 VDPWR.n31 VDPWR 0.076587
R1242 VDPWR.n2 VDPWR 0.076587
R1243 VDPWR.n40 VDPWR 0.0558125
R1244 VDPWR.n34 VDPWR 0.0498421
R1245 VDPWR.n5 VDPWR 0.0498421
R1246 VDPWR.n69 VDPWR.n39 0.0483835
R1247 VDPWR.n107 VDPWR 0.0483723
R1248 VDPWR.n152 VDPWR 0.0483723
R1249 VDPWR VDPWR.n31 0.0465526
R1250 VDPWR VDPWR.n2 0.0465526
R1251 VDPWR.n66 VDPWR 0.0199611
R1252 VDPWR.n83 VDPWR 0.0199611
R1253 VDPWR.n31 VDPWR.n30 0.0168043
R1254 VDPWR.n2 VDPWR.n1 0.0168043
R1255 VDPWR.n68 VDPWR.n40 0.014875
R1256 VDPWR.n125 VDPWR.n124 0.0135682
R1257 VDPWR.n24 VDPWR.n23 0.0135682
R1258 VDPWR.n28 VDPWR 0.0121279
R1259 VDPWR.n35 VDPWR.n34 0.00707895
R1260 VDPWR.n6 VDPWR.n5 0.00707895
R1261 VDPWR.n66 VDPWR.n53 0.00499102
R1262 VDPWR.n83 VDPWR.n70 0.00499102
R1263 VDPWR.n38 VDPWR.n37 0.00340698
R1264 VDPWR.n155 VDPWR.n8 0.00321739
R1265 VDPWR VDPWR.n156 0.00321739
R1266 VDPWR VDPWR.n106 0.00116489
R1267 VDPWR VDPWR.n151 0.00116489
R1268 ua[0].n6 ua[0].n4 2724.21
R1269 ua[0].n9 ua[0].n8 2724.21
R1270 ua[0].n7 ua[0].n6 1018.07
R1271 ua[0].n9 ua[0].n3 1018.07
R1272 ua[0].n12 ua[0].t3 649.886
R1273 ua[0].n0 ua[0].t1 649.692
R1274 ua[0].n5 ua[0].n1 526.307
R1275 ua[0].n5 ua[0].n2 526.307
R1276 ua[0].n10 ua[0].n2 497.486
R1277 ua[0].n11 ua[0].n1 493.762
R1278 ua[0].n6 ua[0].n5 37.0005
R1279 ua[0].n10 ua[0].n9 37.0005
R1280 ua[0].n14 ua[0] 13.435
R1281 ua[0].n4 ua[0].n1 5.78175
R1282 ua[0].n8 ua[0].n2 5.78175
R1283 ua[0].n0 ua[0].t0 4.69622
R1284 ua[0].n4 ua[0].n3 3.61407
R1285 ua[0].n8 ua[0].n7 3.61407
R1286 ua[0].t2 ua[0].n3 2.16152
R1287 ua[0].n7 ua[0].t2 2.16152
R1288 ua[0].n12 ua[0].n11 1.8605
R1289 ua[0].n11 ua[0].n10 1.54533
R1290 ua[0].n14 ua[0].n13 0.9005
R1291 ua[0].n13 ua[0].n0 0.64055
R1292 ua[0].n13 ua[0].n12 0.405262
R1293 ua[0] ua[0].n14 0.0639375
R1294 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t2 669.481
R1295 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t0 669.481
R1296 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t3 218.06
R1297 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t1 218.06
R1298 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t9 211.017
R1299 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t8 208.394
R1300 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t6 208.394
R1301 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t4 207.43
R1302 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t7 207.43
R1303 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t5 207.43
R1304 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t0 649.773
R1305 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t5 649.691
R1306 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.n3 594.383
R1307 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.n4 594.301
R1308 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t6 227.361
R1309 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t8 216.731
R1310 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t13 216.731
R1311 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t14 216.731
R1312 flash_0.x7.neg_mid_b.n0 flash_0.x7.neg_mid_b.t15 105.956
R1313 flash_0.x7.neg_mid_b.n2 flash_0.x7.neg_mid_b 103.529
R1314 flash_0.x7.neg_mid_b.t8 flash_0.x7.neg_mid_b.t7 101.221
R1315 flash_0.x7.neg_mid_b.t13 flash_0.x7.neg_mid_b.t11 101.221
R1316 flash_0.x7.neg_mid_b.t14 flash_0.x7.neg_mid_b.t12 101.221
R1317 flash_0.x7.neg_mid_b.n4 flash_0.x7.neg_mid_b.t4 55.3905
R1318 flash_0.x7.neg_mid_b.n4 flash_0.x7.neg_mid_b.t2 55.3905
R1319 flash_0.x7.neg_mid_b.n3 flash_0.x7.neg_mid_b.t3 55.3905
R1320 flash_0.x7.neg_mid_b.n3 flash_0.x7.neg_mid_b.t1 55.3905
R1321 flash_0.x7.neg_mid_b.n2 flash_0.x7.neg_mid_b.n1 22.3887
R1322 flash_0.x7.neg_mid_b.n1 flash_0.x7.neg_mid_b.t10 8.4355
R1323 flash_0.x7.neg_mid_b.n1 flash_0.x7.neg_mid_b.t9 8.4355
R1324 flash_0.x7.neg_mid_b.n0 flash_0.x7.neg_mid_b 5.14452
R1325 flash_0.x7.neg_mid_b.n0 flash_0.x7.neg_mid_b.n2 2.45104
R1326 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.n0 1.98963
R1327 flash_0.x6.Y flash_0.x6.Y.t0 84.4155
R1328 flash_0.x5.A.n6 flash_0.x5.A.n4 2888.05
R1329 flash_0.x5.A.n9 flash_0.x5.A.n3 2888.05
R1330 flash_0.x5.A.n11 flash_0.x5.A.t3 658.039
R1331 flash_0.x5.A.n8 flash_0.x5.A.n4 509.978
R1332 flash_0.x5.A.n7 flash_0.x5.A.n3 509.978
R1333 flash_0.x5.A.n5 flash_0.x5.A.n2 334.683
R1334 flash_0.x5.A.n10 flash_0.x5.A.n2 334.683
R1335 flash_0.x5.A.n5 flash_0.x5.A.n1 291.084
R1336 flash_0.x5.A.n1 flash_0.x5.A.n10 290.635
R1337 flash_0.x5.A.n0 flash_0.x5.A.t0 215.056
R1338 flash_0.x5.A.n6 flash_0.x5.A.n5 146.25
R1339 flash_0.x5.A.n10 flash_0.x5.A.n9 146.25
R1340 flash_0.x5.A.n7 flash_0.x5.A.n6 114.621
R1341 flash_0.x5.A.n9 flash_0.x5.A.n8 114.621
R1342 flash_0.x5.A flash_0.x5.A.t4 33.6612
R1343 flash_0.x5.A flash_0.x5.A.t5 32.9049
R1344 flash_0.x5.A.n4 flash_0.x5.A.n2 32.5005
R1345 flash_0.x5.A.n3 flash_0.x5.A.n1 32.5005
R1346 flash_0.x5.A.t1 flash_0.x5.A.n7 25.8261
R1347 flash_0.x5.A.n8 flash_0.x5.A.t1 25.8261
R1348 flash_0.x5.A.n0 flash_0.x5.A.t2 17.2847
R1349 flash_0.x5.A flash_0.x5.A.n11 2.49814
R1350 flash_0.x5.A.n0 flash_0.x5.A.n1 1.43573
R1351 flash_0.x5.A.n11 flash_0.x5.A.n0 1.12981
R1352 ui_in[0].n0 ui_in[0].t6 207.43
R1353 ui_in[0].n1 ui_in[0].t14 207.43
R1354 ui_in[0].n2 ui_in[0].t8 207.43
R1355 ui_in[0].n3 ui_in[0].t9 207.43
R1356 ui_in[0].n4 ui_in[0].t0 207.43
R1357 ui_in[0].n5 ui_in[0].t10 207.43
R1358 ui_in[0].n26 ui_in[0].n23 123.867
R1359 ui_in[0].n25 ui_in[0] 50.8126
R1360 ui_in[0].n15 ui_in[0] 50.8126
R1361 ui_in[0] ui_in[0].n1 48.5522
R1362 ui_in[0] ui_in[0].n3 48.5522
R1363 ui_in[0].n6 ui_in[0].n5 47.7953
R1364 ui_in[0].n6 ui_in[0].n2 32.1435
R1365 ui_in[0].n8 ui_in[0] 29.9794
R1366 ui_in[0].n10 ui_in[0] 29.9794
R1367 ui_in[0].n21 ui_in[0] 29.418
R1368 ui_in[0].n18 ui_in[0] 29.418
R1369 ui_in[0].n27 ui_in[0] 26.7297
R1370 ui_in[0].n25 ui_in[0].n24 19.0005
R1371 ui_in[0].n21 ui_in[0].n20 19.0005
R1372 ui_in[0].n18 ui_in[0].n17 19.0005
R1373 ui_in[0].n15 ui_in[0].n14 19.0005
R1374 ui_in[0].n8 ui_in[0].n7 19.0005
R1375 ui_in[0].n10 ui_in[0].n9 19.0005
R1376 ui_in[0] ui_in[0].n0 13.6833
R1377 ui_in[0] ui_in[0].n4 13.6833
R1378 ui_in[0].n20 ui_in[0].t17 12.0505
R1379 ui_in[0].n20 ui_in[0].t15 12.0505
R1380 ui_in[0].n17 ui_in[0].t7 12.0505
R1381 ui_in[0].n17 ui_in[0].t4 12.0505
R1382 ui_in[0].n7 ui_in[0].t16 12.0505
R1383 ui_in[0].n7 ui_in[0].t12 12.0505
R1384 ui_in[0].n9 ui_in[0].t5 12.0505
R1385 ui_in[0].n9 ui_in[0].t2 12.0505
R1386 ui_in[0] ui_in[0].n13 11.4683
R1387 ui_in[0].n24 ui_in[0].t13 8.4355
R1388 ui_in[0].n24 ui_in[0].t11 8.4355
R1389 ui_in[0].n14 ui_in[0].t3 8.4355
R1390 ui_in[0].n14 ui_in[0].t1 8.4355
R1391 ui_in[0] ui_in[0].n26 4.94473
R1392 ui_in[0].n13 ui_in[0].n12 4.5005
R1393 ui_in[0].n13 ui_in[0] 4.0005
R1394 ui_in[0].n2 ui_in[0] 3.75222
R1395 ui_in[0].n1 ui_in[0] 3.75222
R1396 ui_in[0].n0 ui_in[0] 3.75222
R1397 ui_in[0].n5 ui_in[0] 3.75222
R1398 ui_in[0].n4 ui_in[0] 3.75222
R1399 ui_in[0].n3 ui_in[0] 3.75222
R1400 ui_in[0].n11 ui_in[0].n8 2.96269
R1401 ui_in[0].n27 ui_in[0] 2.12895
R1402 ui_in[0].n12 ui_in[0].n6 1.69929
R1403 ui_in[0].n16 ui_in[0].n15 1.59032
R1404 ui_in[0].n22 ui_in[0].n19 1.42722
R1405 ui_in[0].n19 ui_in[0].n18 1.32907
R1406 ui_in[0].n22 ui_in[0].n21 1.32907
R1407 ui_in[0].n26 ui_in[0].n25 1.32907
R1408 ui_in[0].n11 ui_in[0].n10 1.32907
R1409 ui_in[0].n23 ui_in[0].n16 1.29347
R1410 ui_in[0].n12 ui_in[0].n11 0.48697
R1411 ui_in[0].n19 ui_in[0].n16 0.25925
R1412 ui_in[0].n23 ui_in[0].n22 0.25925
R1413 ui_in[0].n13 ui_in[0] 0.0611061
R1414 ui_in[0] ui_in[0].n27 0.02925
R1415 flash_0.x7.VOUT.n8 flash_0.x7.VOUT.n6 2045.32
R1416 flash_0.x7.VOUT.n11 flash_0.x7.VOUT.n5 2045.32
R1417 flash_0.x7.VOUT.n9 flash_0.x7.VOUT.n8 836.909
R1418 flash_0.x7.VOUT.n11 flash_0.x7.VOUT.n10 836.909
R1419 flash_0.x7.VOUT flash_0.x7.VOUT.t6 649.691
R1420 flash_0.x7.VOUT flash_0.x7.VOUT.t9 649.691
R1421 flash_0.x7.VOUT flash_0.x7.VOUT.t14 649.691
R1422 flash_0.x7.VOUT flash_0.x7.VOUT.t8 649.691
R1423 flash_0.x7.VOUT flash_0.x7.VOUT.n2 594.383
R1424 flash_0.x7.VOUT flash_0.x7.VOUT.n13 594.301
R1425 flash_0.x7.VOUT flash_0.x7.VOUT.n14 594.301
R1426 flash_0.x7.VOUT flash_0.x7.VOUT.n3 594.301
R1427 flash_0.x7.VOUT flash_0.x7.VOUT.t1 227.431
R1428 flash_0.x7.VOUT flash_0.x7.VOUT.t2 227.361
R1429 flash_0.x7.VOUT.n6 flash_0.x7.VOUT.n4 195
R1430 flash_0.x7.VOUT.n12 flash_0.x7.VOUT.n11 146.25
R1431 flash_0.x7.VOUT.n8 flash_0.x7.VOUT.n7 146.25
R1432 flash_0.x7.VOUT.n12 flash_0.x7.VOUT.n4 132.894
R1433 flash_0.x7.VOUT.n7 flash_0.x7.VOUT.n4 132.894
R1434 flash_0.x7.VOUT.n9 flash_0.x7.VOUT.n5 105.183
R1435 flash_0.x7.VOUT.n10 flash_0.x7.VOUT.n6 105.183
R1436 flash_0.x7.VOUT.n12 flash_0.x7.VOUT.n1 53.1377
R1437 flash_0.x7.VOUT.n10 flash_0.x7.VOUT.t0 79.7913
R1438 flash_0.x7.VOUT.t0 flash_0.x7.VOUT.n9 79.7913
R1439 flash_0.x7.VOUT.n13 flash_0.x7.VOUT.t7 55.3905
R1440 flash_0.x7.VOUT.n13 flash_0.x7.VOUT.t5 55.3905
R1441 flash_0.x7.VOUT.n14 flash_0.x7.VOUT.t3 55.3905
R1442 flash_0.x7.VOUT.n14 flash_0.x7.VOUT.t4 55.3905
R1443 flash_0.x7.VOUT.n3 flash_0.x7.VOUT.t12 55.3905
R1444 flash_0.x7.VOUT.n3 flash_0.x7.VOUT.t11 55.3905
R1445 flash_0.x7.VOUT.n2 flash_0.x7.VOUT.t10 55.3905
R1446 flash_0.x7.VOUT.n2 flash_0.x7.VOUT.t13 55.3905
R1447 flash_0.x7.VOUT.n7 flash_0.x7.VOUT.n0 52.7987
R1448 flash_0.x7.VOUT flash_0.x7.VOUT.n0 28.5614
R1449 flash_0.x7.VOUT.n0 flash_0.x7.VOUT.n1 0.446827
R1450 flash_0.x7.VOUT.n5 flash_0.x7.VOUT.n1 198.951
R1451 w_7728_24730.t2 w_7728_24730.t0 336.07
R1452 w_7728_24730.t1 w_7728_24730.t2 649.856
R1453 w_7728_24730.t2 w_7728_24730.t3 649.692
R1454 flash_0.x3.clka flash_0.x3.clka.t0 167.038
R1455 flash_0.x3.clka flash_0.x3.clka.t1 87.4292
R1456 flash_0.x3.clkb flash_0.x3.clkb.t0 167.038
R1457 flash_0.x3.clkb flash_0.x3.clkb.t1 87.4292
R1458 flash_0.x4.pos_en_b.n0 flash_0.x4.pos_en_b.t0 669.481
R1459 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.t1 669.481
R1460 flash_0.x4.pos_en_b flash_0.x4.pos_en_b.t3 218.06
R1461 flash_0.x4.pos_en_b flash_0.x4.pos_en_b.t2 218.06
R1462 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.t4 65.4032
R1463 flash_0.x4.pos_en_b.t4 flash_0.x4.pos_en_b 56.2429
R1464 flash_0.x4.pos_en_b.t4 flash_0.x4.pos_en_b 56.2429
R1465 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b 50.8126
R1466 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b 50.8126
R1467 flash_0.x4.pos_en_b flash_0.x4.pos_en_b.n1 29.0914
R1468 flash_0.x4.pos_en_b.n0 flash_0.x4.pos_en_b 29.0914
R1469 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.n0 28.2591
R1470 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.t5 27.4355
R1471 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.t6 27.4355
R1472 ui_in[2].n1 ui_in[2].t1 150.088
R1473 ui_in[2].n0 ui_in[2].t2 33.6007
R1474 ui_in[2].n0 ui_in[2].t0 32.9049
R1475 ui_in[2].n2 ui_in[2] 31.3871
R1476 ui_in[2].n2 ui_in[2].n1 4.55612
R1477 ui_in[2].n1 ui_in[2] 1.9712
R1478 ui_in[2] ui_in[2].n0 0.063
R1479 ui_in[2] ui_in[2].n2 0.047375
R1480 flash_0.x2.clka flash_0.x2.clka.t0 167.038
R1481 flash_0.x2.clka flash_0.x2.clka.t1 87.4292
R1482 flash_0.x7.dcgint.n0 flash_0.x7.dcgint.t4 644.461
R1483 flash_0.x7.dcgint.n5 flash_0.x7.dcgint.t1 640.39
R1484 flash_0.x7.dcgint.n3 flash_0.x7.dcgint.n1 605.365
R1485 flash_0.x7.dcgint.n3 flash_0.x7.dcgint.n2 605.365
R1486 flash_0.x7.dcgint.n4 flash_0.x7.dcgint.t0 477.228
R1487 flash_0.x7.dcgint.t0 flash_0.x7.dcgint.t2 339.594
R1488 flash_0.x7.dcgint.t2 flash_0.x7.dcgint.t6 339.594
R1489 flash_0.x7.dcgint flash_0.x7.dcgint.t11 227.361
R1490 flash_0.x7.dcgint flash_0.x7.dcgint.t10 227.361
R1491 flash_0.x7.dcgint flash_0.x7.dcgint.t9 227.361
R1492 flash_0.x7.dcgint.n4 flash_0.x7.dcgint.n3 69.5657
R1493 flash_0.x7.dcgint.n1 flash_0.x7.dcgint.t3 55.3905
R1494 flash_0.x7.dcgint.n1 flash_0.x7.dcgint.t7 55.3905
R1495 flash_0.x7.dcgint.n2 flash_0.x7.dcgint.t5 55.3905
R1496 flash_0.x7.dcgint.n2 flash_0.x7.dcgint.t8 55.3905
R1497 flash_0.x7.dcgint.n6 flash_0.x7.dcgint.n5 9.3005
R1498 flash_0.x7.dcgint.n5 flash_0.x7.dcgint.n4 8.9605
R1499 flash_0.x7.dcgint flash_0.x7.dcgint.n6 7.52362
R1500 flash_0.x7.dcgint.n6 flash_0.x7.dcgint.n0 1.14684
R1501 flash_0.x7.dcgint.n4 flash_0.x7.dcgint.n0 1.0086
R1502 uo_out[0].n0 uo_out[0].t0 228.901
R1503 uo_out[0].n0 uo_out[0].t1 84.4155
R1504 uo_out[0].n1 uo_out[0] 32.5825
R1505 uo_out[0].n1 uo_out[0].n0 4.88722
R1506 uo_out[0].n0 uo_out[0] 0.063
R1507 uo_out[0] uo_out[0].n1 0.016125
C0 uo_out[0] flash_0.x7.VPRGNEG 3.06829f
C1 flash_0.x7.VPRGPOS flash_0.x4.pos_mid_b 2.26733f
C2 flash_0.x7.neg_en_b ui_in[0] 3.05692f
C3 VAPWR flash_0.x2.clkinb 1.65827f
C4 flash_0.x4.VOUT flash_0.x7.VPRGPOS 1.81318f
C5 flash_0.x2.stage1 flash_0.x2.clka 57.610302f
C6 flash_0.x4.VOUT VDPWR 2.67515f
C7 flash_0.x7.VOUT flash_0.x7.VPRGPOS 4.05693f
C8 VDPWR flash_0.x7.neg_mid 1.38354f
C9 flash_0.x6.Y VDPWR 7.946081f
C10 VDPWR flash_0.x4.neg_en_b 1.82688f
C11 flash_0.x2.clkb flash_0.x2.clka 1.38778f
C12 VAPWR flash_0.x2.stage1 5.931509f
C13 flash_0.x3.stage1 flash_0.x3.clka 57.6093f
C14 flash_0.x3.clka flash_0.x3.clkb 1.38778f
C15 VDPWR flash_0.x7.VOUT 2.37329f
C16 flash_0.x4.neg_mid_b flash_0.x4.neg_mid 1.16207f
C17 flash_0.x7.neg_en_b flash_0.x7.neg_mid 1.5384f
C18 VAPWR flash_0.x3.clka 1.5347f
C19 flash_0.x7.VOUT flash_0.x7.VPRGNEG 1.06096f
C20 flash_0.x3.stage2 flash_0.x7.VPRGPOS 1.93468f
C21 ui_in[2] clk 2.12761f
C22 VDPWR flash_0.x4.neg_mid 1.39258f
C23 VAPWR flash_0.x3.clkina 1.05609f
C24 VDPWR flash_0.x7.neg_mid_b 1.80655f
C25 clk flash_0.x3.stage1 1.05122f
C26 VDPWR flash_0.x4.pos_en_b 1.88599f
C27 flash_0.x7.VPRGNEG flash_0.x7.neg_mid_b 2.18563f
C28 flash_0.x4.neg_mid_b ui_in[1] 1.66762f
C29 flash_0.x3.stage1 flash_0.x3.stage2 5.8896f
C30 flash_0.x3.stage2 flash_0.x3.clkb 59.0307f
C31 clk VAPWR 2.76692f
C32 VAPWR flash_0.x3.stage2 1.42027f
C33 flash_0.x2.stage1 flash_0.x3.clka 4.27357f
C34 flash_0.x2.clka flash_0.x2.stage2 1.79536f
C35 flash_0.x7.VPRGNEG flash_0.x2.stage2 1.79888f
C36 ui_in[2] ui_in[1] 4.33387f
C37 VDPWR ui_in[1] 3.76549f
C38 clk ui_in[0] 4.50971f
C39 VAPWR flash_0.x2.clkina 1.04794f
C40 flash_0.x7.pos_en_b ui_in[1] 2.34386f
C41 flash_0.x3.clkb flash_0.x2.stage2 4.24817f
C42 VAPWR flash_0.x2.stage2 7.897181f
C43 VDPWR flash_0.x4.neg_mid_b 1.91965f
C44 ui_in[0] flash_0.x7.neg_mid_b 1.58977f
C45 clk flash_0.x2.stage1 2.76362f
C46 flash_0.x4.pos_en_b ui_in[0] 2.34221f
C47 flash_0.x7.neg_mid_b flash_0.x7.dcgint 2.14914f
C48 flash_0.x4.neg_mid_b flash_0.x7.VPRGNEG 2.19355f
C49 VDPWR flash_0.x7.VPRGPOS 3.90775f
C50 flash_0.x7.VPRGPOS flash_0.x7.VPRGNEG 1.33754f
C51 flash_0.x3.stage2 flash_0.x3.clka 1.79536f
C52 ui_in[2] VDPWR 3.57578f
C53 VDPWR flash_0.x7.VPRGNEG 13.5121f
C54 VDPWR flash_0.x7.pos_en_b 1.83158f
C55 ui_in[0] ui_in[1] 8.14454f
C56 flash_0.x4.neg_en_b flash_0.x4.neg_mid 1.5384f
C57 flash_0.x4.pos_mid flash_0.x4.pos_mid_b 1.82667f
C58 flash_0.x7.neg_en_b VDPWR 1.68116f
C59 flash_0.x2.stage1 flash_0.x2.stage2 4.80565f
C60 flash_0.x7.neg_mid flash_0.x7.neg_mid_b 1.16207f
C61 flash_0.x5.A flash_0.x7.VPRGPOS 2.9732f
C62 VAPWR flash_0.x7.VPRGNEG 2.20506f
C63 flash_0.x5.A VDPWR 2.1939f
C64 VAPWR flash_0.x3.clkinb 1.66476f
C65 uo_out[0] flash_0.x7.VPRGPOS 2.61882f
C66 flash_0.x2.clkb flash_0.x2.stage2 58.9902f
C67 VAPWR flash_0.x3.stage1 4.90996f
C68 flash_0.x7.pos_mid_b flash_0.x7.VPRGPOS 2.35676f
C69 uo_out[0] ui_in[2] 2.38891f
C70 flash_0.x4.neg_en_b ui_in[1] 3.07359f
C71 flash_0.x7.pos_mid_b flash_0.x7.pos_mid 1.82667f
C72 flash_0.x4.dcgint flash_0.x4.neg_mid_b 2.14914f
C73 VDPWR ui_in[0] 3.61976f
C74 ui_in[0] VGND 23.163868f
C75 ui_in[1] VGND 20.608742f
C76 uo_out[0] VGND 13.615086f
C77 ui_in[2] VGND 15.806785f
C78 clk VGND 25.498615f
C79 ua[0] VGND 35.369205f
C80 VDPWR VGND 0.100366p
C81 VAPWR VGND 43.180836f
C82 flash_0.x7.pos_mid VGND 1.29172f
C83 flash_0.x7.pos_mid_b VGND 3.990245f
C84 flash_0.x4.pos_mid VGND 1.32119f
C85 flash_0.x4.pos_mid_b VGND 4.041469f
C86 flash_0.x6.Y VGND 13.6985f
C87 flash_0.x7.neg_en_b VGND 3.319396f
C88 flash_0.x7.neg_mid_b VGND 4.331881f
C89 flash_0.x7.pos_en_b VGND 7.751863f
C90 flash_0.x4.neg_en_b VGND 3.199904f
C91 flash_0.x4.neg_mid_b VGND 4.866097f
C92 flash_0.x4.pos_en_b VGND 7.775064f
C93 flash_0.x4.VOUT VGND 7.269768f
C94 flash_0.x2.clkb VGND 63.13064f
C95 flash_0.x2.clka VGND 62.52466f
C96 flash_0.x2.clkinb VGND 3.11026f
C97 flash_0.x2.clkina VGND 1.57797f
C98 flash_0.x3.clkb VGND 66.16767f
C99 flash_0.x3.clka VGND 65.171394f
C100 flash_0.x3.clkinb VGND 3.10612f
C101 flash_0.x3.clkina VGND 1.5755f
C102 flash_0.x7.dcgint VGND 3.318307f
C103 flash_0.x4.dcgint VGND 2.996747f
C104 flash_0.x5.A VGND 5.742692f
C105 flash_0.x7.VOUT VGND 12.946657f
C106 flash_0.x7.VPRGNEG VGND 80.182205f
C107 flash_0.x2.stage2 VGND 15.4695f
C108 flash_0.x2.stage1 VGND 18.413f
C109 flash_0.x7.VPRGPOS VGND 0.148816p
C110 flash_0.x3.stage2 VGND 24.3058f
C111 flash_0.x3.stage1 VGND 23.173801f
C112 uo_out[0].n1 VGND 3.39873f
C113 ui_in[2].n1 VGND 1.125f
C114 ui_in[2].n2 VGND 4.50156f
C115 w_7728_24730.t0 VGND 6.5007f
C116 w_7728_24730.t2 VGND 6.37557f
C117 flash_0.x7.VOUT.n0 VGND 2.13265f
C118 ui_in[0].n13 VGND 1.02386f
C119 ui_in[0].n27 VGND 3.82492f
C120 ua[0].n14 VGND 1.92631f
C121 VDPWR.n39 VGND 12.558001f
C122 VDPWR.n46 VGND 1.02977f
C123 VDPWR.t53 VGND 1.65275f
C124 VDPWR.n49 VGND 1.02977f
C125 VDPWR.n69 VGND 1.05184f
C126 VDPWR.n84 VGND 1.56105f
C127 ui_in[1].n27 VGND 4.6267f
C128 clk.n2 VGND 1.74152f
C129 clk.n3 VGND 4.1318f
C130 VAPWR.n123 VGND 1.0575f
C131 VAPWR.n125 VGND 7.2806f
C132 VAPWR.n126 VGND 40.983803f
C133 flash_0.x7.VPRGPOS.n17 VGND 2.01105f
.ends

