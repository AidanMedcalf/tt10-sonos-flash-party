* NGSPICE file created from charge_pump_neg_nmos.ext - technology: sky130A

.subckt charge_pump_neg_nmos clk VOUT VAPWR VGND
X0 clkina clkinb VAPWR.t5 VAPWR.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X1 clkinb clk.t0 VGND.t1 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X2 stage1 stage1 VGND.t9 stage1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 stage2 stage2 stage1 stage2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 clkb clkinb VGND.t5 VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X5 clkb clkinb VAPWR.t3 VAPWR.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X6 VOUT VGND.t6 sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X7 VOUT.t2 VOUT.t0 stage2 VOUT.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X8 clkinb clk.t1 VAPWR.t1 VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X9 clkina clkinb VGND.t3 VGND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X10 clka clkina VGND.t8 VGND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X11 clka clkina VAPWR.t6 VAPWR.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X12 clkb stage2 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X13 clka stage1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
R0 VAPWR.n6 VAPWR.n5 2332.91
R1 VAPWR.n7 VAPWR.n6 2332.91
R2 VAPWR.n8 VAPWR.n7 2332.91
R3 VAPWR.n8 VAPWR.n5 2332.91
R4 VAPWR.n6 VAPWR.n0 29.5749
R5 VAPWR.n9 VAPWR.n4 1551.32
R6 VAPWR.n9 VAPWR.n2 15.7169
R7 VAPWR.n0 VAPWR.t5 649.99
R8 VAPWR.n0 VAPWR.t1 649.765
R9 VAPWR.t0 VAPWR.t4 487.901
R10 VAPWR.n1 VAPWR.n0 38.8984
R11 VAPWR.t0 VAPWR.n0 355.545
R12 VAPWR.n2 VAPWR.n5 25.2299
R13 VAPWR.n3 VAPWR.n0 96.11
R14 VAPWR VAPWR.n0 96.096
R15 VAPWR VAPWR.n0 95.7547
R16 VAPWR.n0 VAPWR.t3 167.41
R17 VAPWR.n0 VAPWR.t6 167.251
R18 VAPWR.n1 VAPWR.t2 2.91292
R19 VAPWR.t4 VAPWR.n1 28.7038
R20 VAPWR.n0 VAPWR.n2 16.641
R21 VAPWR.n9 VAPWR.n8 14.2313
R22 VAPWR.n0 VAPWR.n4 12.116
R23 VAPWR.n7 VAPWR.n4 12.3338
R24 clk clk.t1 54.3383
R25 clk clk.t0 53.1307
R26 VGND.n3 VGND.n7 17010.2
R27 VGND.n8 VGND.n7 17010.2
R28 VGND.n13 VGND.n12 9438.3
R29 VGND.n12 VGND.n11 5607.68
R30 VGND.n12 VGND.n5 4686.84
R31 VGND.n13 VGND.t6 193.419
R32 VGND.t6 VGND.n1 47.2327
R33 VGND.n6 VGND.n5 3370.76
R34 VGND.n11 VGND.n9 2547.06
R35 VGND.n9 VGND.n6 2166.87
R36 VGND.n7 VGND.n6 1472.95
R37 VGND.t6 VGND.n2 7.29093
R38 VGND.n11 VGND.n10 957.745
R39 VGND.t4 VGND.t7 838.864
R40 VGND.t2 VGND.t0 838.864
R41 VGND.n10 VGND.t4 530.34
R42 VGND.n13 VGND.t0 530.34
R43 VGND.t7 VGND.n1 419.433
R44 VGND.n1 VGND.t2 419.433
R45 VGND.t6 VGND.t3 227.643
R46 VGND.t6 VGND.t1 227.398
R47 VGND.n10 VGND.t6 195.087
R48 VGND.t6 VGND.t8 82.9558
R49 VGND.n0 VGND.t9 78.1972
R50 VGND.n0 VGND.n14 33.1299
R51 VGND.n4 VGND.n3 9.28621
R52 VGND.n3 VGND.n5 9.28621
R53 VGND.n8 VGND.t6 9.28621
R54 VGND.n9 VGND.n8 9.28621
R55 VGND.n2 VGND.n4 8.15439
R56 VGND.t6 VGND.n0 6.2055
R57 VGND.n4 VGND 5.97887
R58 VGND.t5 VGND.t6 83.1878
R59 VGND.n2 VGND.n7 27.0289
R60 VGND.t6 VGND 12.3552
R61 VOUT.n1 VOUT.n3 808.657
R62 VOUT.n4 VOUT.n2 837.184
R63 VOUT VOUT.t0 113.356
R64 VOUT.n4 VOUT.n1 200.702
R65 VOUT.n3 VOUT.n2 198.256
R66 VOUT VOUT.t2 82.8472
R67 VOUT VOUT.n2 10.785
R68 VOUT.t1 VOUT.n3 66.988
R69 VOUT.n4 VOUT.t1 66.988
R70 VOUT VOUT.n0 17.2678
R71 VOUT.n1 VOUT 12.7784
C0 VAPWR stage1 3.79319f
C1 VAPWR stage2 7.8754f
C2 VAPWR VOUT 2.15626f
C3 stage2 clkb 58.9902f
C4 clka stage1 57.615f
C5 stage2 stage1 4.80565f
C6 VOUT VGND 74.50468f
C7 VAPWR VGND 29.73482f
C8 clkb VGND 4.7031f
C9 clka VGND 5.27941f
C10 clkinb VGND 3.10612f
C11 stage2 VGND 17.2767f
C12 stage1 VGND 16.4132f
C13 VAPWR.n0 VGND 9.66749f
.ends

