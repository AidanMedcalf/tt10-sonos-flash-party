* NGSPICE file created from tt_um_sonos_flash_party.ext - technology: sky130A

.subckt tt_um_sonos_flash_party clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VDPWR VGND VAPWR
X0 flash_0.x7.VPRGNEG VGND.t42 sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X1 flash_0.x7.VPRGPOS.t28 flash_0.x7.pos_mid_b.t3 flash_0.x7.vintp flash_0.x7.VPRGPOS.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X2 flash_0.x2.clkb.t1 flash_0.x2.clkinb VAPWR.t15 VAPWR.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X3 flash_0.x7.VPRGPOS.t30 flash_0.x7.pos_mid flash_0.x7.pos_mid_b.t2 flash_0.x7.VPRGPOS.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X4 flash_0.x3.clkinb clk.t0 VAPWR.t12 VAPWR.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X5 flash_0.x7.VPRGPOS.t29 flash_0.x4.pos_mid flash_0.x4.pos_mid_b.t2 flash_0.x7.VPRGPOS.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X6 VGND.t66 ui_in[1].t0 flash_0.x4.neg_en_b.t1 VGND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X7 flash_0.x4.dcgint.t8 flash_0.x4.neg_mid_b.t7 flash_0.x4.VOUT.t8 flash_0.x4.dcgint.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X8 flash_0.x7.pos_mid_b.t1 ui_in[1].t1 VGND.t39 VGND.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X9 flash_0.x7.pos_mid flash_0.x7.pos_en_b.t4 VGND.t69 VGND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X10 VDPWR.t44 ui_in[1].t2 flash_0.x4.neg_mid VDPWR.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X11 ua[0].t1 VGND.t40 VGND.t41 ua[0].t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=10
X12 VDPWR.t48 flash_0.x7.neg_en_b.t4 flash_0.x7.neg_mid_b.t5 VDPWR.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X13 VDPWR.t28 flash_0.x7.neg_en_b.t5 flash_0.x7.neg_mid_b.t4 VDPWR.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X14 flash_0.x5.A.t0 flash_0.x6.Y VDPWR.t46 VDPWR.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
X15 flash_0.x7.vintp flash_0.x7.pos_mid_b.t4 flash_0.x7.VPRGPOS.t27 flash_0.x7.VPRGPOS.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X16 flash_0.x7.neg_mid ui_in[0].t0 VDPWR.t3 VDPWR.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X17 flash_0.x4.neg_mid_b.t6 flash_0.x4.neg_mid flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=1
X18 flash_0.x2.clkina flash_0.x2.clkinb VAPWR.t14 VAPWR.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X19 flash_0.x4.neg_mid_b.t2 flash_0.x4.neg_en_b.t4 VDPWR.t23 VDPWR.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X20 flash_0.x7.pos_mid_b.t0 ui_in[1].t3 VGND.t24 VGND.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X21 flash_0.x7.pos_mid flash_0.x7.pos_en_b.t4 VGND.t68 VGND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X22 flash_0.x4.dcgint.t7 flash_0.x4.neg_mid_b.t8 flash_0.x4.VOUT.t12 flash_0.x4.dcgint.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X23 a_9352_28387# flash_0.x4.VOUT.t14 a_7463_28281# flash_0.x7.VOUT.t14 sky130_fd_bs_flash__special_sonosfet_star ad=0.13725 pd=1.51 as=0.13725 ps=1.51 w=0.45 l=0.22
X24 VGND.t17 ui_in[1].t4 flash_0.x7.pos_mid_b VGND.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X25 VGND.t1 ui_in[0].t1 flash_0.x4.pos_mid_b VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X26 flash_0.x7.VPRGNEG flash_0.x4.neg_mid_b.t9 flash_0.x4.neg_mid flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.145 ps=1.58 w=0.5 l=1
X27 flash_0.x4.vintp VDPWR flash_0.x4.VOUT.t6 flash_0.x7.VPRGPOS.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X28 VDPWR.t43 ui_in[1].t5 flash_0.x4.neg_en_b.t2 VDPWR.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X29 flash_0.x4.VOUT.t0 VDPWR.t58 a_16296_28578# flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X30 VDPWR.t52 flash_0.x7.neg_en_b.t6 flash_0.x7.neg_mid_b.t3 VDPWR.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X31 w_7728_24730.t3 ua[0].t2 ua[0].t3 w_7728_24730.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
X32 flash_0.x3.stage1 VAPWR.t8 VAPWR.t10 VAPWR.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X33 flash_0.x4.VOUT.t5 VDPWR flash_0.x4.vintp flash_0.x7.VPRGPOS.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X34 flash_0.x7.neg_en_b.t0 ui_in[0].t2 VGND.t25 VGND.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X35 flash_0.x7.pos_en_b.t2 ui_in[1].t6 VGND.t3 VGND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X36 VGND.t11 ui_in[1].t7 flash_0.x7.pos_mid_b VGND.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X37 flash_0.x3.clka.t1 flash_0.x3.clkina VAPWR.t16 VAPWR.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X38 VGND.t27 ui_in[0].t3 flash_0.x4.pos_mid_b VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X39 flash_0.x3.clkb.t0 flash_0.x3.clkinb VGND.t46 VGND.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X40 flash_0.x4.vintp flash_0.x4.pos_mid_b.t3 flash_0.x7.VPRGPOS.t12 flash_0.x7.VPRGPOS.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X41 flash_0.x4.VOUT.t7 VDPWR.t59 a_16296_28578# flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X42 flash_0.x4.dcgint.t11 flash_0.x4.pos_en_b.t4 VGND.t64 VGND.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X43 flash_0.x7.VPRGPOS.t3 flash_0.x4.pos_mid_b.t4 flash_0.x4.vintp flash_0.x7.VPRGPOS.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X44 flash_0.x6.Y.t0 ui_in[2].t0 VGND.t48 VGND.t47 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X45 flash_0.x7.VOUT.t7 VDPWR flash_0.x7.vintp flash_0.x7.VPRGPOS.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X46 flash_0.x2.clka.t0 flash_0.x2.clkina VGND.t38 VGND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X47 flash_0.x3.clkb flash_0.x3.stage2 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X48 VGND.t67 ui_in[1].t8 flash_0.x7.pos_en_b.t1 VGND.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X49 VGND.t16 ui_in[0].t4 flash_0.x4.pos_en_b.t3 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X50 VDPWR.t21 flash_0.x4.neg_en_b.t5 flash_0.x4.neg_mid_b.t3 VDPWR.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X51 flash_0.x7.neg_en_b.t2 ui_in[0].t5 VDPWR.t50 VDPWR.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=3
X52 flash_0.x7.pos_en_b.t3 ui_in[1].t9 VDPWR.t41 VDPWR.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X53 flash_0.x4.dcgint.t10 flash_0.x4.pos_en_b.t4 VGND.t62 VGND.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X54 VDPWR.t39 ui_in[1].t10 flash_0.x4.neg_mid VDPWR.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X55 a_16296_28578# flash_0.x4.neg_mid_b.t10 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X56 flash_0.x4.neg_mid_b.t5 flash_0.x4.neg_en_b.t6 VDPWR.t19 VDPWR.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X57 flash_0.x7.VPRGPOS.t26 flash_0.x7.pos_mid_b.t5 flash_0.x7.vintp flash_0.x7.VPRGPOS.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X58 flash_0.x7.neg_mid ui_in[0].t6 VDPWR.t10 VDPWR.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X59 flash_0.x4.neg_mid_b.t0 flash_0.x4.neg_en_b.t7 VDPWR.t17 VDPWR.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X60 flash_0.x4.dcgint.t5 flash_0.x4.neg_mid_b.t11 flash_0.x4.VOUT.t13 flash_0.x4.dcgint.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X61 flash_0.x7.VPRGPOS.t9 w_7728_24730.t0 w_7728_24730.t1 flash_0.x7.VPRGPOS.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
X62 VDPWR.t38 ui_in[1].t11 flash_0.x7.pos_en_b.t0 VDPWR.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X63 flash_0.x3.clkinb clk.t1 VGND.t19 VGND.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X64 VDPWR.t30 ui_in[0].t7 flash_0.x4.pos_en_b.t1 VDPWR.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X65 flash_0.x2.clkina flash_0.x2.clkinb VGND.t52 VGND.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X66 flash_0.x3.clka flash_0.x3.stage1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X67 a_16296_28578# flash_0.x4.neg_mid_b.t10 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X68 flash_0.x4.dcgint.t9 flash_0.x4.pos_en_b.t4 VGND.t60 VGND.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X69 flash_0.x4.VOUT.t9 flash_0.x4.neg_mid_b.t12 flash_0.x4.dcgint.t4 flash_0.x4.dcgint.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X70 flash_0.x4.dcgint.t3 flash_0.x4.neg_mid_b.t13 flash_0.x4.VOUT.t11 flash_0.x4.dcgint.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X71 flash_0.x4.vintp VDPWR flash_0.x4.VOUT.t4 flash_0.x7.VPRGPOS.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X72 a_7463_28281# ui_in[2].t1 VGND.t22 VGND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X73 flash_0.x7.neg_mid ui_in[0].t8 VDPWR.t11 VDPWR.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X74 flash_0.x7.dcgint.t11 flash_0.x7.neg_mid_b.t7 flash_0.x7.VOUT.t11 flash_0.x7.dcgint.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X75 VDPWR.t57 ui_in[0].t9 flash_0.x7.neg_mid VDPWR.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X76 uo_out[0].t0 flash_0.x5.A.t4 VDPWR.t5 VDPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X77 VDPWR.t56 ui_in[0].t10 flash_0.x7.neg_mid VDPWR.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X78 flash_0.x4.VOUT.t3 VDPWR flash_0.x4.vintp flash_0.x7.VPRGPOS.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X79 flash_0.x3.stage2 flash_0.x3.stage1 flash_0.x3.stage1 flash_0.x3.stage1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X80 flash_0.x2.clkinb clk.t2 VAPWR.t1 VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X81 flash_0.x4.VOUT.t10 flash_0.x4.neg_mid_b.t14 flash_0.x4.dcgint.t1 flash_0.x4.dcgint.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X82 flash_0.x7.neg_mid_b.t6 flash_0.x7.neg_mid flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=1
X83 flash_0.x4.vintp flash_0.x4.pos_mid_b.t5 flash_0.x7.VPRGPOS.t31 flash_0.x7.VPRGPOS.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X84 VGND.t55 flash_0.x7.pos_en_b.t5 flash_0.x7.pos_mid VGND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X85 flash_0.x7.dcgint.t10 flash_0.x7.neg_mid_b.t8 flash_0.x7.VOUT.t12 flash_0.x7.dcgint.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X86 flash_0.x3.clkb.t1 flash_0.x3.clkinb VAPWR.t7 VAPWR.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X87 flash_0.x7.vintp VDPWR flash_0.x7.VOUT.t6 flash_0.x7.VPRGPOS.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X88 flash_0.x7.VOUT.t1 VDPWR.t60 a_20416_28577# flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X89 flash_0.x4.vintp VDPWR flash_0.x4.VOUT.t2 flash_0.x7.VPRGPOS.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X90 flash_0.x7.VPRGPOS.t1 flash_0.x4.pos_mid_b.t6 flash_0.x4.vintp flash_0.x7.VPRGPOS.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X91 flash_0.x2.clkb flash_0.x2.stage2 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X92 flash_0.x2.stage1 flash_0.x2.stage1 VGND.t20 flash_0.x2.stage1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X93 flash_0.x7.VPRGPOS.t10 flash_0.x3.stage2 flash_0.x3.stage2 flash_0.x3.stage2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X94 VGND.t54 flash_0.x7.pos_en_b.t5 flash_0.x7.pos_mid VGND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X95 flash_0.x4.pos_mid_b.t1 ui_in[0].t11 VGND.t26 VGND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X96 flash_0.x4.pos_mid flash_0.x4.pos_en_b.t5 VGND.t31 VGND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X97 flash_0.x2.clkb.t0 flash_0.x2.clkinb VGND.t50 VGND.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X98 flash_0.x3.clkina flash_0.x3.clkinb VAPWR.t5 VAPWR.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X99 flash_0.x7.vintp flash_0.x7.pos_mid_b.t6 flash_0.x7.VPRGPOS.t25 flash_0.x7.VPRGPOS.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X100 VDPWR.t15 flash_0.x4.neg_en_b.t8 flash_0.x4.neg_mid_b.t1 VDPWR.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X101 flash_0.x7.VOUT.t0 VDPWR.t61 a_20416_28577# flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X102 flash_0.x4.vintp flash_0.x4.pos_mid_b.t7 flash_0.x7.VPRGPOS.t7 flash_0.x7.VPRGPOS.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X103 flash_0.x7.dcgint.t2 flash_0.x7.pos_en_b.t6 VGND.t9 VGND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X104 a_20416_28577# flash_0.x7.neg_mid_b.t9 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X105 flash_0.x2.clka.t1 flash_0.x2.clkina VAPWR.t3 VAPWR.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X106 VGND.t56 ui_in[0].t12 flash_0.x7.neg_en_b.t3 VGND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X107 flash_0.x7.neg_mid_b.t2 flash_0.x7.neg_en_b.t7 VDPWR.t8 VDPWR.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X108 flash_0.x4.pos_mid_b.t0 ui_in[0].t13 VGND.t13 VGND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X109 flash_0.x4.neg_mid ui_in[1].t12 VDPWR.t36 VDPWR.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X110 flash_0.x4.pos_mid flash_0.x4.pos_en_b.t5 VGND.t30 VGND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X111 VDPWR.t35 ui_in[1].t13 flash_0.x4.neg_mid VDPWR.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X112 flash_0.x2.clka flash_0.x2.stage1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X113 flash_0.x7.VPRGPOS VGND.t70 sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X114 VDPWR.t13 flash_0.x4.neg_en_b.t9 flash_0.x4.neg_mid_b.t4 VDPWR.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X115 flash_0.x7.dcgint.t1 flash_0.x7.pos_en_b.t6 VGND.t7 VGND.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X116 a_20416_28577# flash_0.x7.neg_mid_b.t10 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X117 flash_0.x7.VOUT.t9 flash_0.x7.neg_mid_b.t11 flash_0.x7.dcgint.t8 flash_0.x7.dcgint.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X118 VDPWR.t55 ui_in[0].t14 flash_0.x7.neg_mid VDPWR.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X119 flash_0.x7.neg_mid_b.t1 flash_0.x7.neg_en_b.t8 VDPWR.t24 VDPWR.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X120 flash_0.x4.neg_en_b.t0 ui_in[1].t14 VGND.t65 VGND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X121 flash_0.x4.pos_en_b.t2 ui_in[0].t15 VGND.t29 VGND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X122 flash_0.x4.neg_mid ui_in[1].t15 VDPWR.t34 VDPWR.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X123 VDPWR.t26 ui_in[0].t16 flash_0.x7.neg_en_b.t1 VDPWR.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X124 flash_0.x7.dcgint.t7 flash_0.x7.neg_mid_b.t12 flash_0.x7.VOUT.t8 flash_0.x7.dcgint.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X125 flash_0.x2.clkinb clk.t3 VGND.t36 VGND.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X126 flash_0.x7.VOUT.t10 flash_0.x7.neg_mid_b.t13 flash_0.x7.dcgint.t6 flash_0.x7.dcgint.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X127 flash_0.x4.VOUT.t1 VDPWR flash_0.x4.vintp flash_0.x7.VPRGPOS.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X128 flash_0.x7.dcgint.t0 flash_0.x7.pos_en_b.t6 VGND.t5 VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X129 flash_0.x3.clka.t0 flash_0.x3.clkina VGND.t58 VGND.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X130 flash_0.x5.A.t3 flash_0.x5.A.t1 a_9352_28387# flash_0.x5.A.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.5
X131 flash_0.x7.dcgint.t4 flash_0.x7.neg_mid_b.t14 flash_0.x7.VOUT.t13 flash_0.x7.dcgint.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X132 flash_0.x7.neg_mid_b.t0 flash_0.x7.neg_en_b.t9 VDPWR.t7 VDPWR.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X133 flash_0.x7.vintp VDPWR flash_0.x7.VOUT.t5 flash_0.x7.VPRGPOS.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X134 flash_0.x4.neg_en_b.t3 ui_in[1].t16 VDPWR.t33 VDPWR.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=3
X135 flash_0.x4.pos_en_b.t0 ui_in[0].t17 VDPWR.t1 VDPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X136 VGND.t34 flash_0.x4.pos_en_b.t6 flash_0.x4.pos_mid VGND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X137 flash_0.x7.VPRGNEG flash_0.x7.neg_mid_b.t15 flash_0.x7.neg_mid flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.145 ps=1.58 w=0.5 l=1
X138 flash_0.x7.VOUT.t4 VDPWR flash_0.x7.vintp flash_0.x7.VPRGPOS.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X139 flash_0.x2.stage2 flash_0.x2.stage2 flash_0.x2.stage1 flash_0.x2.stage2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X140 flash_0.x7.VPRGPOS.t32 flash_0.x4.pos_mid_b.t8 flash_0.x4.vintp flash_0.x7.VPRGPOS.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X141 flash_0.x4.neg_mid ui_in[1].t17 VDPWR.t31 VDPWR.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X142 flash_0.x7.vintp flash_0.x7.pos_mid_b.t7 flash_0.x7.VPRGPOS.t24 flash_0.x7.VPRGPOS.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X143 flash_0.x7.VOUT.t3 VDPWR flash_0.x7.vintp flash_0.x7.VPRGPOS.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X144 flash_0.x7.VPRGPOS.t23 flash_0.x7.pos_mid_b flash_0.x7.pos_mid flash_0.x7.VPRGPOS.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X145 flash_0.x7.VPRGPOS.t5 flash_0.x4.pos_mid_b flash_0.x4.pos_mid flash_0.x7.VPRGPOS.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X146 VGND.t33 flash_0.x4.pos_en_b.t6 flash_0.x4.pos_mid VGND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X147 uo_out[0].t1 flash_0.x5.A.t5 VGND.t15 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X148 flash_0.x3.clkina flash_0.x3.clkinb VGND.t44 VGND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X149 flash_0.x7.vintp VDPWR flash_0.x7.VOUT.t2 flash_0.x7.VPRGPOS.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X150 flash_0.x7.VPRGPOS.t21 flash_0.x7.pos_mid_b.t8 flash_0.x7.vintp flash_0.x7.VPRGPOS.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X151 flash_0.x6.Y ui_in[2].t2 VDPWR.t54 VDPWR.t53 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X152 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG flash_0.x2.stage2 flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
R0 VGND.t59 VGND.n121 1.77808e+07
R1 VGND.n211 VGND.n210 1.32662e+07
R2 VGND.n121 VGND.t4 9.06413e+06
R3 VGND.n211 VGND.n24 7.77048e+06
R4 VGND.n138 VGND.n129 136400
R5 VGND.n152 VGND.n118 77206.1
R6 VGND.n178 VGND.n63 55379.3
R7 VGND.n140 VGND.n139 41452.9
R8 VGND.n136 VGND.n135 28158.7
R9 VGND.n82 VGND.n67 26564
R10 VGND.n143 VGND.n129 26182
R11 VGND.n82 VGND.n81 19464
R12 VGND.n139 VGND.n138 18707.2
R13 VGND.n177 VGND.n176 17794
R14 VGND.n212 VGND.n22 17579
R15 VGND.n45 VGND.n41 17010.2
R16 VGND.n52 VGND.n41 17010.2
R17 VGND.n189 VGND.n56 17010.2
R18 VGND.n180 VGND.n56 17010.2
R19 VGND.n148 VGND.n129 16052.9
R20 VGND.n136 VGND.n22 15944.1
R21 VGND.n176 VGND.n82 15655.2
R22 VGND.n158 VGND.n118 15267.5
R23 VGND.n178 VGND.n177 13983.9
R24 VGND.n177 VGND.n64 12678.4
R25 VGND.n138 VGND.n137 11203.8
R26 VGND.n213 VGND.n212 8682.25
R27 VGND.n158 VGND.n157 8288.46
R28 VGND.n71 VGND.n22 7672.91
R29 VGND.n128 VGND.t63 6465.71
R30 VGND.n137 VGND.n118 5878.85
R31 VGND.n211 VGND.n23 5801.34
R32 VGND.n58 VGND.n55 5607.68
R33 VGND.n43 VGND.n40 5607.68
R34 VGND.n40 VGND.n23 5607.68
R35 VGND.n62 VGND.n55 5607.68
R36 VGND.n120 VGND.n119 5067.26
R37 VGND.n141 VGND.n140 4557.14
R38 VGND.t53 VGND.t2 4288.33
R39 VGND.t2 VGND.t10 4288.33
R40 VGND.t32 VGND.t28 4288.33
R41 VGND.t28 VGND.t0 4288.33
R42 VGND.n174 VGND.n83 3957.38
R43 VGND.n174 VGND.n84 3957.38
R44 VGND.n133 VGND.n84 3957.38
R45 VGND.n133 VGND.n83 3957.38
R46 VGND.n72 VGND.n68 3957.38
R47 VGND.n72 VGND.n69 3957.38
R48 VGND.n80 VGND.n69 3957.38
R49 VGND.n80 VGND.n68 3957.38
R50 VGND.n209 VGND.n25 3790.36
R51 VGND.n60 VGND.n25 3790.36
R52 VGND.n195 VGND.n194 3790.36
R53 VGND.n194 VGND.n38 3790.36
R54 VGND.n151 VGND.t23 3495.43
R55 VGND.n142 VGND.t12 3495.43
R56 VGND.n81 VGND.t47 3200.66
R57 VGND.n71 VGND.t47 3200.66
R58 VGND.n152 VGND.n151 2827
R59 VGND.n143 VGND.n142 2827
R60 VGND.n43 VGND.n39 2736.73
R61 VGND.n150 VGND.n148 2648.22
R62 VGND.n139 VGND.n135 2546
R63 VGND.t10 VGND.n150 2345.18
R64 VGND.t0 VGND.n141 2345.18
R65 VGND.n178 VGND.n62 2341.85
R66 VGND.n157 VGND.t23 2331.85
R67 VGND.n63 VGND.n58 2309.11
R68 VGND.n54 VGND.n53 2233.78
R69 VGND.n137 VGND.n136 2176.84
R70 VGND.n212 VGND.n211 1977.24
R71 VGND.n214 VGND.n20 1900.12
R72 VGND.n214 VGND.n21 1900.12
R73 VGND.n66 VGND.n21 1900.12
R74 VGND.n66 VGND.n20 1900.12
R75 VGND.n191 VGND.n190 1830.35
R76 VGND.t12 VGND.n128 1820.3
R77 VGND.n140 VGND.n64 1788.04
R78 VGND.n135 VGND.n134 1768.36
R79 VGND.n44 VGND.n23 1501.04
R80 VGND.n54 VGND.n39 1195.35
R81 VGND.n176 VGND.n175 1151.51
R82 VGND.n51 VGND.n42 1139.95
R83 VGND.n46 VGND.n42 1139.95
R84 VGND.n188 VGND.n57 1139.95
R85 VGND.n181 VGND.n57 1139.95
R86 VGND.t8 VGND.n158 1094.37
R87 VGND.n134 VGND.t14 1089.55
R88 VGND.n175 VGND.t14 1089.55
R89 VGND.n120 VGND.n54 931.699
R90 VGND.n62 VGND.n61 883.615
R91 VGND.n151 VGND.t53 792.894
R92 VGND.n142 VGND.t32 792.894
R93 VGND.t49 VGND.t37 757.616
R94 VGND.n67 VGND.t21 660
R95 VGND.n213 VGND.t21 660
R96 VGND.n179 VGND.n58 657.409
R97 VGND.n15 VGND.t41 650.87
R98 VGND.t51 VGND.t35 597.753
R99 VGND.n147 VGND.n144 535.718
R100 VGND.n156 VGND.n153 535.718
R101 VGND.n121 VGND.n120 522.082
R102 VGND.t63 VGND.t61 487.856
R103 VGND.n61 VGND.t49 478.974
R104 VGND.t57 VGND.t45 470.42
R105 VGND.n208 VGND.n207 437.836
R106 VGND.n207 VGND.n27 437.836
R107 VGND.n197 VGND.n37 437.836
R108 VGND.n197 VGND.n196 437.836
R109 VGND.n210 VGND.t35 424.973
R110 VGND.n44 VGND.n43 417.728
R111 VGND.n191 VGND.n54 402.44
R112 VGND.t37 VGND.n59 378.808
R113 VGND.n59 VGND.t51 378.808
R114 VGND.t43 VGND.t18 350.719
R115 VGND.n127 VGND.t59 304.329
R116 VGND.t45 VGND.n192 297.404
R117 VGND.n132 VGND.n131 257.13
R118 VGND.n132 VGND.n86 257.13
R119 VGND.n79 VGND.n70 257.13
R120 VGND.n79 VGND.n78 257.13
R121 VGND.n193 VGND.t57 235.209
R122 VGND.n163 VGND.t5 230.898
R123 VGND.n161 VGND.t7 230.898
R124 VGND.n162 VGND.t9 230.898
R125 VGND.n125 VGND.t60 230.898
R126 VGND.n122 VGND.t62 230.898
R127 VGND.n123 VGND.t64 230.898
R128 VGND.n131 VGND.n85 229.272
R129 VGND.n172 VGND.n86 229.272
R130 VGND.n74 VGND.n70 229.272
R131 VGND.n78 VGND.n77 229.272
R132 VGND.n199 VGND.t44 227.643
R133 VGND.n205 VGND.t52 227.643
R134 VGND.n26 VGND.t36 227.398
R135 VGND.n34 VGND.t19 227.398
R136 VGND.n193 VGND.t43 222.901
R137 VGND.n215 VGND.n19 221.742
R138 VGND.n65 VGND.n19 221.742
R139 VGND.n65 VGND.n18 221.742
R140 VGND.t18 VGND.n24 221.728
R141 VGND.n144 VGND.n143 188.038
R142 VGND.n153 VGND.n152 188.038
R143 VGND.t61 VGND.n127 183.528
R144 VGND.n148 VGND.n147 180.132
R145 VGND.n157 VGND.n156 180.132
R146 VGND.t6 VGND.t8 157.787
R147 VGND.n216 VGND.n18 152.194
R148 VGND.n150 VGND.n149 152.111
R149 VGND.n141 VGND.n130 152.111
R150 VGND.n135 VGND.n64 147.569
R151 VGND.n20 VGND.n18 146.25
R152 VGND.t21 VGND.n20 146.25
R153 VGND.n21 VGND.n19 146.25
R154 VGND.t21 VGND.n21 146.25
R155 VGND.n133 VGND.n132 117.001
R156 VGND.n134 VGND.n133 117.001
R157 VGND.n174 VGND.n173 117.001
R158 VGND.n175 VGND.n174 117.001
R159 VGND.n80 VGND.n79 117.001
R160 VGND.n81 VGND.n80 117.001
R161 VGND.n73 VGND.n72 117.001
R162 VGND.n72 VGND.n71 117.001
R163 VGND.n192 VGND.n191 107.427
R164 VGND.n53 VGND.n40 102.35
R165 VGND.n190 VGND.n55 102.35
R166 VGND.n159 VGND.t4 98.4295
R167 VGND.n60 VGND.n27 97.5005
R168 VGND.n61 VGND.n60 97.5005
R169 VGND.n209 VGND.n208 97.5005
R170 VGND.n210 VGND.n209 97.5005
R171 VGND.n38 VGND.n37 97.5005
R172 VGND.n192 VGND.n38 97.5005
R173 VGND.n196 VGND.n195 97.5005
R174 VGND.n195 VGND.n24 97.5005
R175 VGND.n115 VGND.n114 97.1505
R176 VGND.n108 VGND.n107 97.1505
R177 VGND.n111 VGND.n110 97.1505
R178 VGND.n104 VGND.n103 97.1505
R179 VGND.n113 VGND.n112 97.1505
R180 VGND.n106 VGND.n105 97.1505
R181 VGND.n99 VGND.n98 97.1505
R182 VGND.n92 VGND.n91 97.1505
R183 VGND.n95 VGND.n94 97.1505
R184 VGND.n88 VGND.n87 97.1505
R185 VGND.n97 VGND.n96 97.1505
R186 VGND.n90 VGND.n89 97.1505
R187 VGND.n119 VGND.n63 95.855
R188 VGND.n114 VGND.t3 95.7605
R189 VGND.n114 VGND.t67 95.7605
R190 VGND.n107 VGND.t25 95.7605
R191 VGND.n107 VGND.t56 95.7605
R192 VGND.n110 VGND.t68 95.7605
R193 VGND.n110 VGND.t11 95.7605
R194 VGND.n103 VGND.t24 95.7605
R195 VGND.n103 VGND.t54 95.7605
R196 VGND.n112 VGND.t69 95.7605
R197 VGND.n112 VGND.t17 95.7605
R198 VGND.n105 VGND.t39 95.7605
R199 VGND.n105 VGND.t55 95.7605
R200 VGND.n98 VGND.t29 95.7605
R201 VGND.n98 VGND.t16 95.7605
R202 VGND.n91 VGND.t65 95.7605
R203 VGND.n91 VGND.t66 95.7605
R204 VGND.n94 VGND.t30 95.7605
R205 VGND.n94 VGND.t27 95.7605
R206 VGND.n87 VGND.t13 95.7605
R207 VGND.n87 VGND.t33 95.7605
R208 VGND.n96 VGND.t31 95.7605
R209 VGND.n96 VGND.t1 95.7605
R210 VGND.n89 VGND.t26 95.7605
R211 VGND.n89 VGND.t34 95.7605
R212 VGND.n170 VGND.t15 83.754
R213 VGND.n76 VGND.t48 83.7172
R214 VGND.n36 VGND.t46 83.1807
R215 VGND.n28 VGND.t50 83.1807
R216 VGND.n35 VGND.t58 82.9558
R217 VGND.n29 VGND.t38 82.9558
R218 VGND.n30 VGND.t20 82.8472
R219 VGND.n160 VGND.n159 73.7068
R220 VGND.n127 VGND.n126 73.7068
R221 VGND.n66 VGND.n65 65.0005
R222 VGND.n67 VGND.n66 65.0005
R223 VGND.n215 VGND.n214 65.0005
R224 VGND.n214 VGND.n213 65.0005
R225 VGND.n159 VGND.t6 59.3584
R226 VGND.n216 VGND.n215 56.9466
R227 VGND.n131 VGND.n83 53.1823
R228 VGND.n83 VGND.t14 53.1823
R229 VGND.n86 VGND.n84 53.1823
R230 VGND.n84 VGND.t14 53.1823
R231 VGND.n70 VGND.n68 53.1823
R232 VGND.n68 VGND.t47 53.1823
R233 VGND.n78 VGND.n69 53.1823
R234 VGND.n69 VGND.t47 53.1823
R235 VGND.n217 VGND.t22 41.2645
R236 VGND.n173 VGND.n85 27.8593
R237 VGND.n173 VGND.n172 27.8593
R238 VGND.n74 VGND.n73 27.8593
R239 VGND.n77 VGND.n73 27.8593
R240 VGND.n57 VGND.n56 26.5914
R241 VGND.n119 VGND.n56 26.5914
R242 VGND.n42 VGND.n41 26.5914
R243 VGND.n41 VGND.n39 26.5914
R244 VGND.n207 VGND.n25 24.3755
R245 VGND.n59 VGND.n25 24.3755
R246 VGND.n197 VGND.n194 24.3755
R247 VGND.n194 VGND.n193 24.3755
R248 VGND.n179 VGND.n178 20.4593
R249 VGND.n75 VGND.n74 9.35514
R250 VGND.n77 VGND 9.33194
R251 VGND.n172 VGND.n171 9.3005
R252 VGND.n171 VGND.n85 9.3005
R253 VGND.n46 VGND.n45 9.28621
R254 VGND.n45 VGND.n44 9.28621
R255 VGND.n189 VGND.n188 9.28621
R256 VGND.n190 VGND.n189 9.28621
R257 VGND.n52 VGND.n51 9.28621
R258 VGND.n53 VGND.n52 9.28621
R259 VGND.n181 VGND.n180 9.28621
R260 VGND.n180 VGND.n179 9.28621
R261 VGND.n219 VGND.n16 8.39735
R262 VGND.n48 VGND.n47 8.21246
R263 VGND.n187 VGND.n186 8.21246
R264 VGND.n49 VGND.n48 7.33652
R265 VGND.n186 VGND.n185 7.33652
R266 VGND.n149 VGND.n117 6.24424
R267 VGND.n130 VGND.n101 6.24424
R268 VGND.n47 VGND 5.82387
R269 VGND.n187 VGND 5.82387
R270 VGND.n218 VGND.n217 5.18907
R271 VGND.n50 VGND 5.15194
R272 VGND.n182 VGND 5.15194
R273 VGND.n170 VGND.n169 5.15155
R274 VGND.n15 VGND.t40 4.756
R275 VGND.n124 VGND.n123 4.5005
R276 VGND.n124 VGND.n122 4.5005
R277 VGND.n125 VGND.n124 4.5005
R278 VGND.n164 VGND.n162 4.5005
R279 VGND.n164 VGND.n161 4.5005
R280 VGND.n164 VGND.n163 4.5005
R281 VGND.n33 VGND.n32 4.12801
R282 VGND.n184 VGND.n183 4.12801
R283 VGND.n150 VGND.n128 4.11265
R284 VGND.n146 VGND.n145 3.83474
R285 VGND.n155 VGND.n154 3.83474
R286 VGND.n202 VGND 3.81988
R287 VGND.n221 VGND 3.32011
R288 VGND.n37 VGND.n36 3.31952
R289 VGND.n28 VGND.n27 3.31952
R290 VGND.n201 VGND.n33 3.218
R291 VGND.n16 VGND.n15 3.20171
R292 VGND.n166 VGND.n165 3.12737
R293 VGND.n168 VGND.n167 3.00925
R294 uio_oe[7] VGND.n221 2.60868
R295 VGND.n217 VGND.n216 2.3255
R296 VGND.n109 VGND.n106 2.2505
R297 VGND.n116 VGND.n113 2.2505
R298 VGND.n109 VGND.n104 2.2505
R299 VGND.n116 VGND.n111 2.2505
R300 VGND.n109 VGND.n108 2.2505
R301 VGND.n116 VGND.n115 2.2505
R302 VGND.n93 VGND.n90 2.2505
R303 VGND.n100 VGND.n97 2.2505
R304 VGND.n93 VGND.n88 2.2505
R305 VGND.n100 VGND.n95 2.2505
R306 VGND.n93 VGND.n92 2.2505
R307 VGND.n100 VGND.n99 2.2505
R308 VGND.n126 VGND.n125 2.04916
R309 VGND.n163 VGND.n160 2.04916
R310 VGND.n169 VGND.n168 2.00487
R311 VGND.n184 VGND.n31 1.913
R312 VGND.n145 VGND.n144 1.8605
R313 VGND.n147 VGND.n146 1.8605
R314 VGND.n156 VGND.n155 1.8605
R315 VGND.n154 VGND.n153 1.8605
R316 VGND.n169 VGND.n17 1.74613
R317 VGND.n31 VGND.n30 1.5555
R318 VGND.n208 VGND.n26 1.5505
R319 VGND.n196 VGND.n34 1.5505
R320 VGND.n166 VGND.n117 1.31425
R321 VGND.n203 VGND.n31 1.3055
R322 VGND.n168 VGND.n101 1.248
R323 VGND.n218 VGND.n17 1.188
R324 VGND.n202 VGND.n17 1.1555
R325 VGND.n36 VGND.n35 0.879043
R326 VGND.n29 VGND.n28 0.879043
R327 VGND.n221 VGND.n220 0.751794
R328 VGND.n219 VGND.n218 0.525188
R329 VGND.n204 VGND.n203 0.501003
R330 VGND.n201 VGND.n200 0.501003
R331 VGND.n48 VGND.n42 0.443357
R332 VGND.n186 VGND.n57 0.443357
R333 VGND.n207 VGND.n206 0.404848
R334 VGND.n198 VGND.n197 0.404848
R335 VGND.n116 VGND.n109 0.378453
R336 VGND.n100 VGND.n93 0.378453
R337 VGND.n145 VGND 0.321152
R338 VGND.n154 VGND 0.321152
R339 VGND.n165 VGND.n160 0.285933
R340 VGND.n126 VGND.n102 0.28175
R341 VGND.n146 VGND 0.280391
R342 VGND.n155 VGND 0.280391
R343 VGND.n167 VGND.n166 0.27425
R344 VGND.n167 VGND.n102 0.236484
R345 VGND.n206 VGND.n205 0.221088
R346 VGND.n199 VGND.n198 0.221088
R347 VGND.n205 VGND 0.214961
R348 VGND VGND.n199 0.214961
R349 VGND.n124 VGND 0.204732
R350 VGND VGND.n164 0.204732
R351 VGND VGND.n202 0.177375
R352 VGND.n75 VGND.n16 0.168469
R353 VGND.n220 VGND.n219 0.166437
R354 VGND.n0 uo_out[1] 0.16627
R355 VGND.n1 uo_out[2] 0.16627
R356 VGND.n2 uo_out[3] 0.16627
R357 VGND.n3 uo_out[4] 0.16627
R358 VGND.n4 uo_out[5] 0.16627
R359 VGND.n5 uo_out[6] 0.16627
R360 VGND.n6 uo_out[7] 0.16627
R361 VGND.n7 uio_out[0] 0.16627
R362 VGND.n8 uio_out[1] 0.16627
R363 VGND.n9 uio_out[2] 0.16627
R364 VGND.n10 uio_out[3] 0.16627
R365 VGND.n11 uio_out[4] 0.16627
R366 VGND.n12 uio_out[5] 0.16627
R367 VGND.n13 uio_out[6] 0.16627
R368 VGND.n14 uio_out[7] 0.16627
R369 uio_oe[0] VGND.n228 0.16627
R370 uio_oe[1] VGND.n227 0.16627
R371 uio_oe[2] VGND.n226 0.16627
R372 uio_oe[3] VGND.n225 0.16627
R373 uio_oe[4] VGND.n224 0.16627
R374 uio_oe[5] VGND.n223 0.16627
R375 uio_oe[6] VGND.n222 0.16627
R376 VGND.n149 VGND 0.157483
R377 VGND.n130 VGND 0.157483
R378 VGND.n50 VGND.n49 0.15675
R379 VGND.n185 VGND.n182 0.15675
R380 VGND.n47 VGND.n46 0.1555
R381 VGND.n51 VGND.n50 0.1555
R382 VGND.n188 VGND.n187 0.1555
R383 VGND.n182 VGND.n181 0.1555
R384 VGND.n115 VGND 0.102773
R385 VGND.n108 VGND 0.102773
R386 VGND.n111 VGND 0.102773
R387 VGND.n104 VGND 0.102773
R388 VGND.n113 VGND 0.102773
R389 VGND.n106 VGND 0.102773
R390 VGND.n99 VGND 0.102773
R391 VGND.n92 VGND 0.102773
R392 VGND.n95 VGND 0.102773
R393 VGND.n88 VGND 0.102773
R394 VGND.n97 VGND 0.102773
R395 VGND.n90 VGND 0.102773
R396 VGND.n204 VGND.n26 0.0904491
R397 VGND.n200 VGND.n34 0.0904491
R398 VGND VGND.n204 0.0659475
R399 VGND.n200 VGND 0.0659475
R400 VGND.n49 VGND.n33 0.0657174
R401 VGND.n185 VGND.n184 0.0657174
R402 VGND.n220 VGND 0.062375
R403 VGND.n30 VGND 0.0609396
R404 VGND VGND.n201 0.05925
R405 VGND.n203 VGND 0.05925
R406 VGND.n161 VGND 0.0544773
R407 VGND.n162 VGND 0.0544773
R408 VGND.n122 VGND 0.0544773
R409 VGND.n123 VGND 0.0544773
R410 VGND.n125 VGND 0.048
R411 VGND.n163 VGND 0.048
R412 VGND.n171 VGND.n170 0.034875
R413 VGND.n183 VGND.t42 0.0314016
R414 VGND.n32 VGND.t70 0.0314016
R415 VGND VGND.n102 0.0312579
R416 VGND.n0 uo_out[2] 0.0302667
R417 VGND.n1 uo_out[3] 0.0302667
R418 VGND.n2 uo_out[4] 0.0302667
R419 VGND.n3 uo_out[5] 0.0302667
R420 VGND.n4 uo_out[6] 0.0302667
R421 VGND.n5 uo_out[7] 0.0302667
R422 VGND.n6 uio_out[0] 0.0302667
R423 VGND.n7 uio_out[1] 0.0302667
R424 VGND.n8 uio_out[2] 0.0302667
R425 VGND.n9 uio_out[3] 0.0302667
R426 VGND.n10 uio_out[4] 0.0302667
R427 VGND.n11 uio_out[5] 0.0302667
R428 VGND.n12 uio_out[6] 0.0302667
R429 VGND.n13 uio_out[7] 0.0302667
R430 VGND.n14 uio_oe[0] 0.0302667
R431 VGND.n228 uio_oe[1] 0.0302667
R432 VGND.n227 uio_oe[2] 0.0302667
R433 VGND.n226 uio_oe[3] 0.0302667
R434 VGND.n225 uio_oe[4] 0.0302667
R435 VGND.n224 uio_oe[5] 0.0302667
R436 VGND.n223 uio_oe[6] 0.0302667
R437 VGND.n222 uio_oe[7] 0.0302667
R438 VGND.n165 VGND 0.0270748
R439 VGND VGND.n76 0.0244521
R440 VGND.n206 VGND.n29 0.0194951
R441 VGND.n198 VGND.n35 0.0194951
R442 VGND.n117 VGND.n116 0.0182165
R443 VGND.n101 VGND.n100 0.0182165
R444 uo_out[2] VGND.n0 0.010027
R445 uo_out[3] VGND.n1 0.010027
R446 uo_out[4] VGND.n2 0.010027
R447 uo_out[5] VGND.n3 0.010027
R448 uo_out[6] VGND.n4 0.010027
R449 uo_out[7] VGND.n5 0.010027
R450 uio_out[0] VGND.n6 0.010027
R451 uio_out[1] VGND.n7 0.010027
R452 uio_out[2] VGND.n8 0.010027
R453 uio_out[3] VGND.n9 0.010027
R454 uio_out[4] VGND.n10 0.010027
R455 uio_out[5] VGND.n11 0.010027
R456 uio_out[6] VGND.n12 0.010027
R457 uio_out[7] VGND.n13 0.010027
R458 uio_oe[0] VGND.n14 0.010027
R459 VGND.n228 uio_oe[1] 0.010027
R460 VGND.n227 uio_oe[2] 0.010027
R461 VGND.n226 uio_oe[3] 0.010027
R462 VGND.n225 uio_oe[4] 0.010027
R463 VGND.n224 uio_oe[5] 0.010027
R464 VGND.n223 uio_oe[6] 0.010027
R465 VGND.n222 uio_oe[7] 0.010027
R466 VGND.n171 VGND 0.008625
R467 VGND.n76 VGND.n75 0.0012485
R468 VGND.n183 VGND 0.000981102
R469 VGND.n32 VGND 0.000981102
R470 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t2 649.691
R471 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t0 227.442
R472 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t1 227.361
R473 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t7 216.731
R474 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t8 216.731
R475 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t6 216.731
R476 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t3 216.731
R477 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t4 216.731
R478 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t5 216.731
R479 flash_0.x7.VPRGPOS.n6 flash_0.x7.VPRGPOS.n4 4689.72
R480 flash_0.x7.VPRGPOS.n9 flash_0.x7.VPRGPOS.n8 4689.72
R481 flash_0.x7.VPRGPOS.n7 flash_0.x7.VPRGPOS.n6 1828.1
R482 flash_0.x7.VPRGPOS.n9 flash_0.x7.VPRGPOS.n3 1828.1
R483 flash_0.x7.VPRGPOS.n5 flash_0.x7.VPRGPOS.n1 902.777
R484 flash_0.x7.VPRGPOS.n5 flash_0.x7.VPRGPOS.n2 902.777
R485 flash_0.x7.VPRGPOS.n10 flash_0.x7.VPRGPOS.n2 880.232
R486 flash_0.x7.VPRGPOS.n11 flash_0.x7.VPRGPOS.n1 874.658
R487 flash_0.x7.VPRGPOS.t16 flash_0.x7.VPRGPOS.t22 809.375
R488 flash_0.x7.VPRGPOS.t19 flash_0.x7.VPRGPOS.t4 809.375
R489 flash_0.x7.VPRGPOS.n12 flash_0.x7.VPRGPOS.t9 649.856
R490 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t32 649.715
R491 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t26 649.715
R492 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t30 649.691
R493 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t23 649.691
R494 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t29 649.691
R495 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t5 649.691
R496 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t31 649.691
R497 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t24 649.691
R498 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n14 594.301
R499 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n13 594.301
R500 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n18 594.301
R501 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n19 594.301
R502 flash_0.x7.VPRGPOS.t13 flash_0.x7.VPRGPOS.t20 246.875
R503 flash_0.x7.VPRGPOS.t14 flash_0.x7.VPRGPOS.t13 246.875
R504 flash_0.x7.VPRGPOS.t18 flash_0.x7.VPRGPOS.t14 246.875
R505 flash_0.x7.VPRGPOS.t15 flash_0.x7.VPRGPOS.t18 246.875
R506 flash_0.x7.VPRGPOS.t6 flash_0.x7.VPRGPOS.t17 246.875
R507 flash_0.x7.VPRGPOS.t2 flash_0.x7.VPRGPOS.t6 246.875
R508 flash_0.x7.VPRGPOS.t11 flash_0.x7.VPRGPOS.t2 246.875
R509 flash_0.x7.VPRGPOS.t0 flash_0.x7.VPRGPOS.t11 246.875
R510 flash_0.x7.VPRGPOS.n0 flash_0.x7.VPRGPOS.t15 237.5
R511 flash_0.x7.VPRGPOS.n15 flash_0.x7.VPRGPOS.t0 237.5
R512 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t10 82.8472
R513 flash_0.x7.VPRGPOS.n14 flash_0.x7.VPRGPOS.t12 55.3905
R514 flash_0.x7.VPRGPOS.n14 flash_0.x7.VPRGPOS.t1 55.3905
R515 flash_0.x7.VPRGPOS.n13 flash_0.x7.VPRGPOS.t7 55.3905
R516 flash_0.x7.VPRGPOS.n13 flash_0.x7.VPRGPOS.t3 55.3905
R517 flash_0.x7.VPRGPOS.n18 flash_0.x7.VPRGPOS.t25 55.3905
R518 flash_0.x7.VPRGPOS.n18 flash_0.x7.VPRGPOS.t21 55.3905
R519 flash_0.x7.VPRGPOS.n19 flash_0.x7.VPRGPOS.t27 55.3905
R520 flash_0.x7.VPRGPOS.n19 flash_0.x7.VPRGPOS.t28 55.3905
R521 flash_0.x7.VPRGPOS.n6 flash_0.x7.VPRGPOS.n5 37.0005
R522 flash_0.x7.VPRGPOS.n10 flash_0.x7.VPRGPOS.n9 37.0005
R523 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n0 16.1367
R524 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n15 16.1367
R525 flash_0.x7.VPRGPOS.n17 flash_0.x7.VPRGPOS 13.9898
R526 flash_0.x7.VPRGPOS.n0 flash_0.x7.VPRGPOS.t16 9.3755
R527 flash_0.x7.VPRGPOS.n15 flash_0.x7.VPRGPOS.t19 9.3755
R528 flash_0.x7.VPRGPOS.n4 flash_0.x7.VPRGPOS.n1 3.03329
R529 flash_0.x7.VPRGPOS.n8 flash_0.x7.VPRGPOS.n2 3.03329
R530 flash_0.x7.VPRGPOS.n16 flash_0.x7.VPRGPOS 2.77904
R531 flash_0.x7.VPRGPOS.n11 flash_0.x7.VPRGPOS.n10 2.70819
R532 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n17 2.54902
R533 flash_0.x7.VPRGPOS.n12 flash_0.x7.VPRGPOS.n11 1.8605
R534 flash_0.x7.VPRGPOS.n4 flash_0.x7.VPRGPOS.n3 1.85038
R535 flash_0.x7.VPRGPOS.n8 flash_0.x7.VPRGPOS.n7 1.85038
R536 flash_0.x7.VPRGPOS.n16 flash_0.x7.VPRGPOS.n12 1.79707
R537 flash_0.x7.VPRGPOS.n17 flash_0.x7.VPRGPOS.n16 1.40849
R538 flash_0.x7.VPRGPOS.t8 flash_0.x7.VPRGPOS.n3 1.18321
R539 flash_0.x7.VPRGPOS.n7 flash_0.x7.VPRGPOS.t8 1.18321
R540 VAPWR.n62 VAPWR.n4 2380.24
R541 VAPWR.n114 VAPWR.n73 2380.24
R542 VAPWR.n64 VAPWR.n4 2376.31
R543 VAPWR.n116 VAPWR.n73 2376.31
R544 VAPWR.n44 VAPWR.n42 2332.91
R545 VAPWR.n45 VAPWR.n44 2332.91
R546 VAPWR.n46 VAPWR.n45 2332.91
R547 VAPWR.n46 VAPWR.n42 2332.91
R548 VAPWR.n27 VAPWR.n25 2332.91
R549 VAPWR.n28 VAPWR.n27 2332.91
R550 VAPWR.n29 VAPWR.n28 2332.91
R551 VAPWR.n29 VAPWR.n25 2332.91
R552 VAPWR.n13 VAPWR.n12 2332.91
R553 VAPWR.n13 VAPWR.n11 2332.91
R554 VAPWR.n93 VAPWR.n92 2332.91
R555 VAPWR.n93 VAPWR.n91 2332.91
R556 VAPWR.n87 VAPWR.n83 1577.4
R557 VAPWR.n84 VAPWR.n81 1577.4
R558 VAPWR.n47 VAPWR.n38 1551.32
R559 VAPWR.n43 VAPWR.n38 1551.32
R560 VAPWR.n26 VAPWR.n24 1551.32
R561 VAPWR.n26 VAPWR.n21 1551.32
R562 VAPWR.n30 VAPWR.n21 1551.32
R563 VAPWR.n30 VAPWR.n24 1551.32
R564 VAPWR.n47 VAPWR.n41 1538.26
R565 VAPWR.n43 VAPWR.n41 1538.26
R566 VAPWR.n58 VAPWR.n7 1516.38
R567 VAPWR.n58 VAPWR.n6 1516.38
R568 VAPWR.n110 VAPWR.n76 1516.38
R569 VAPWR.n110 VAPWR.n75 1516.38
R570 VAPWR.n14 VAPWR.n7 1514.88
R571 VAPWR.n14 VAPWR.n6 1514.88
R572 VAPWR.n94 VAPWR.n76 1514.88
R573 VAPWR.n94 VAPWR.n75 1514.88
R574 VAPWR.n12 VAPWR.n5 1046.2
R575 VAPWR.n11 VAPWR.n5 1046.2
R576 VAPWR.n92 VAPWR.n74 1046.2
R577 VAPWR.n91 VAPWR.n74 1046.2
R578 VAPWR.n85 VAPWR.n84 722.497
R579 VAPWR.n87 VAPWR.n86 722.497
R580 VAPWR.n0 VAPWR.t14 649.99
R581 VAPWR.n121 VAPWR.t5 649.99
R582 VAPWR.n1 VAPWR.t1 649.765
R583 VAPWR.n71 VAPWR.t12 649.765
R584 VAPWR.t0 VAPWR.t13 487.901
R585 VAPWR.t11 VAPWR.t4 487.901
R586 VAPWR.n66 VAPWR.n3 460.425
R587 VAPWR.n118 VAPWR.n72 460.425
R588 VAPWR.n66 VAPWR.n65 459.671
R589 VAPWR.n118 VAPWR.n117 459.671
R590 VAPWR.n40 VAPWR.n37 386.635
R591 VAPWR.n48 VAPWR.n40 386.635
R592 VAPWR.n49 VAPWR.n37 386.635
R593 VAPWR.n23 VAPWR.n20 386.635
R594 VAPWR.n31 VAPWR.n23 386.635
R595 VAPWR.n32 VAPWR.n20 386.635
R596 VAPWR.n15 VAPWR.n8 386.635
R597 VAPWR.n15 VAPWR.n9 386.635
R598 VAPWR.n57 VAPWR.n8 386.635
R599 VAPWR.n57 VAPWR.n9 386.635
R600 VAPWR.n95 VAPWR.n77 386.635
R601 VAPWR.n95 VAPWR.n78 386.635
R602 VAPWR.n109 VAPWR.n78 386.635
R603 VAPWR.n109 VAPWR.n77 386.635
R604 VAPWR.n64 VAPWR.t0 331.582
R605 VAPWR.n116 VAPWR.t11 331.582
R606 VAPWR.n61 VAPWR.n60 251.28
R607 VAPWR.n113 VAPWR.n112 251.28
R608 VAPWR.t8 VAPWR 236.188
R609 VAPWR.n97 VAPWR.t8 236.011
R610 VAPWR.n49 VAPWR 195.012
R611 VAPWR.n32 VAPWR 195.012
R612 VAPWR VAPWR.n48 191.625
R613 VAPWR VAPWR.n31 191.625
R614 VAPWR.n106 VAPWR.n82 184.847
R615 VAPWR.n107 VAPWR.n106 184.847
R616 VAPWR.n107 VAPWR.n80 184.847
R617 VAPWR.n82 VAPWR.n80 184.847
R618 VAPWR.n59 VAPWR.n5 172.655
R619 VAPWR.n111 VAPWR.n74 172.655
R620 VAPWR.n55 VAPWR.t15 167.41
R621 VAPWR.n79 VAPWR.t7 167.41
R622 VAPWR.n120 VAPWR.t16 167.251
R623 VAPWR.n68 VAPWR.t3 167.141
R624 VAPWR.n60 VAPWR.n59 160.495
R625 VAPWR.n112 VAPWR.n111 160.495
R626 VAPWR.n107 VAPWR.n81 146.25
R627 VAPWR.n83 VAPWR.n82 146.25
R628 VAPWR.n106 VAPWR.n87 97.5005
R629 VAPWR.n84 VAPWR.n80 97.5005
R630 VAPWR.n105 VAPWR.t10 82.8472
R631 VAPWR.t13 VAPWR.t2 81.0585
R632 VAPWR.t4 VAPWR.t6 81.0585
R633 VAPWR.n85 VAPWR.n83 72.5386
R634 VAPWR.n86 VAPWR.n81 72.5386
R635 VAPWR.n86 VAPWR.t9 66.988
R636 VAPWR.t9 VAPWR.n85 66.988
R637 VAPWR.n63 VAPWR.n61 34.0449
R638 VAPWR.n115 VAPWR.n113 34.0449
R639 VAPWR.n62 VAPWR.n3 23.1255
R640 VAPWR.n63 VAPWR.n62 23.1255
R641 VAPWR.n65 VAPWR.n64 23.1255
R642 VAPWR.n114 VAPWR.n72 23.1255
R643 VAPWR.n115 VAPWR.n114 23.1255
R644 VAPWR.n117 VAPWR.n116 23.1255
R645 VAPWR.t13 VAPWR.n61 21.1116
R646 VAPWR.t4 VAPWR.n113 21.1116
R647 VAPWR.n43 VAPWR.n37 14.2313
R648 VAPWR.n44 VAPWR.n43 14.2313
R649 VAPWR.n48 VAPWR.n47 14.2313
R650 VAPWR.n47 VAPWR.n46 14.2313
R651 VAPWR.n26 VAPWR.n20 14.2313
R652 VAPWR.n27 VAPWR.n26 14.2313
R653 VAPWR.n31 VAPWR.n30 14.2313
R654 VAPWR.n30 VAPWR.n29 14.2313
R655 VAPWR.n15 VAPWR.n14 14.2313
R656 VAPWR.n14 VAPWR.n13 14.2313
R657 VAPWR.n58 VAPWR.n57 14.2313
R658 VAPWR.n59 VAPWR.n58 14.2313
R659 VAPWR.n95 VAPWR.n94 14.2313
R660 VAPWR.n94 VAPWR.n93 14.2313
R661 VAPWR.n110 VAPWR.n109 14.2313
R662 VAPWR.n111 VAPWR.n110 14.2313
R663 VAPWR.n41 VAPWR.n40 12.3338
R664 VAPWR.n42 VAPWR.n41 12.3338
R665 VAPWR.n49 VAPWR.n38 12.3338
R666 VAPWR.n45 VAPWR.n38 12.3338
R667 VAPWR.n24 VAPWR.n23 12.3338
R668 VAPWR.n25 VAPWR.n24 12.3338
R669 VAPWR.n32 VAPWR.n21 12.3338
R670 VAPWR.n28 VAPWR.n21 12.3338
R671 VAPWR.n8 VAPWR.n6 12.3338
R672 VAPWR.n11 VAPWR.n6 12.3338
R673 VAPWR.n9 VAPWR.n7 12.3338
R674 VAPWR.n12 VAPWR.n7 12.3338
R675 VAPWR.n78 VAPWR.n76 12.3338
R676 VAPWR.n92 VAPWR.n76 12.3338
R677 VAPWR.n77 VAPWR.n75 12.3338
R678 VAPWR.n91 VAPWR.n75 12.3338
R679 VAPWR.n66 VAPWR.n4 7.70883
R680 VAPWR.n60 VAPWR.n4 7.70883
R681 VAPWR.n118 VAPWR.n73 7.70883
R682 VAPWR.n112 VAPWR.n73 7.70883
R683 VAPWR.n125 VAPWR 4.11654
R684 VAPWR.n126 VAPWR 4.06671
R685 VAPWR.n123 VAPWR 3.16715
R686 VAPWR.n123 VAPWR 3.13288
R687 VAPWR.n39 VAPWR.n35 2.77496
R688 VAPWR.n39 VAPWR.n36 2.77496
R689 VAPWR.n50 VAPWR.n36 2.77496
R690 VAPWR.n22 VAPWR.n18 2.77496
R691 VAPWR.n22 VAPWR.n19 2.77496
R692 VAPWR.n33 VAPWR.n19 2.77496
R693 VAPWR.n16 VAPWR.n10 2.77496
R694 VAPWR.n17 VAPWR.n16 2.77496
R695 VAPWR.n98 VAPWR.n82 2.3255
R696 VAPWR.n108 VAPWR.n107 2.3255
R697 VAPWR.n54 VAPWR.n3 2.1216
R698 VAPWR.n89 VAPWR.n72 2.09672
R699 VAPWR.n52 VAPWR.n34 1.88425
R700 VAPWR.n106 VAPWR.n105 1.5505
R701 VAPWR.n10 VAPWR 1.40267
R702 VAPWR.n53 VAPWR.n52 1.37675
R703 VAPWR.n96 VAPWR.n95 1.32345
R704 VAPWR.n53 VAPWR.n17 1.23691
R705 VAPWR.n51 VAPWR.n50 1.22254
R706 VAPWR.n34 VAPWR.n33 1.22254
R707 VAPWR.n65 VAPWR.n1 1.163
R708 VAPWR.n117 VAPWR.n71 1.163
R709 VAPWR.n124 VAPWR.n123 1.07737
R710 VAPWR.n51 VAPWR.n35 0.894522
R711 VAPWR.n34 VAPWR.n18 0.894522
R712 VAPWR.n48 VAPWR.n35 0.845955
R713 VAPWR.n37 VAPWR.n36 0.845955
R714 VAPWR.n31 VAPWR.n18 0.845955
R715 VAPWR.n20 VAPWR.n19 0.845955
R716 VAPWR.n16 VAPWR.n15 0.845955
R717 VAPWR.n57 VAPWR.n56 0.845955
R718 VAPWR.n109 VAPWR.n108 0.845955
R719 VAPWR.t2 VAPWR.n63 0.81108
R720 VAPWR.t6 VAPWR.n115 0.81108
R721 VAPWR.n104 VAPWR.n103 0.797375
R722 VAPWR.n40 VAPWR.n39 0.664786
R723 VAPWR.n50 VAPWR.n49 0.664786
R724 VAPWR.n23 VAPWR.n22 0.664786
R725 VAPWR.n33 VAPWR.n32 0.664786
R726 VAPWR.n10 VAPWR.n9 0.664786
R727 VAPWR.n17 VAPWR.n8 0.664786
R728 VAPWR.n101 VAPWR.n78 0.664786
R729 VAPWR.n90 VAPWR.n77 0.664786
R730 VAPWR.n52 VAPWR.n51 0.5005
R731 VAPWR VAPWR.n126 0.491143
R732 VAPWR VAPWR.n88 0.490083
R733 VAPWR.n70 VAPWR.n1 0.448327
R734 VAPWR.n67 VAPWR.n66 0.404848
R735 VAPWR.n119 VAPWR.n118 0.404848
R736 VAPWR.n98 VAPWR.n97 0.3455
R737 VAPWR.n68 VAPWR.n0 0.313
R738 VAPWR.n125 VAPWR.n124 0.2968
R739 VAPWR.n103 VAPWR.n102 0.203625
R740 VAPWR.n96 VAPWR.n90 0.198256
R741 VAPWR.n70 VAPWR.n0 0.188
R742 VAPWR.n55 VAPWR.n54 0.179291
R743 VAPWR.n99 VAPWR.n98 0.163
R744 VAPWR.n56 VAPWR.n2 0.157262
R745 VAPWR.n119 VAPWR 0.152375
R746 VAPWR.n69 VAPWR.n68 0.143
R747 VAPWR.n101 VAPWR.n100 0.14175
R748 VAPWR.n70 VAPWR.n69 0.140949
R749 VAPWR VAPWR.n2 0.136533
R750 VAPWR.n104 VAPWR.n88 0.130708
R751 VAPWR VAPWR.n121 0.123855
R752 VAPWR VAPWR.n70 0.105837
R753 VAPWR.n90 VAPWR.n89 0.0951602
R754 VAPWR.n103 VAPWR.n101 0.0905
R755 VAPWR.n89 VAPWR.n79 0.0695895
R756 VAPWR.n121 VAPWR.n120 0.0690307
R757 VAPWR.n124 VAPWR 0.0651875
R758 VAPWR.n67 VAPWR.n2 0.062375
R759 VAPWR.n105 VAPWR 0.0568725
R760 VAPWR.n100 VAPWR.n99 0.0544216
R761 VAPWR.n122 VAPWR.n71 0.0533274
R762 VAPWR.n97 VAPWR 0.043
R763 VAPWR.n100 VAPWR 0.0364477
R764 VAPWR.n105 VAPWR 0.0364477
R765 VAPWR.n120 VAPWR.n119 0.033625
R766 VAPWR.n99 VAPWR.n96 0.0305
R767 VAPWR.n102 VAPWR 0.029875
R768 VAPWR.n56 VAPWR.n55 0.0297008
R769 VAPWR VAPWR.n122 0.0235263
R770 VAPWR VAPWR.n88 0.0212668
R771 VAPWR.n88 VAPWR 0.01927
R772 VAPWR VAPWR.n104 0.0184739
R773 VAPWR.n102 VAPWR 0.0152764
R774 VAPWR.n108 VAPWR.n79 0.0118818
R775 VAPWR.n108 VAPWR 0.00728914
R776 VAPWR.n122 VAPWR 0.00488596
R777 VAPWR.n54 VAPWR.n53 0.00425
R778 VAPWR.n126 VAPWR.n125 0.0033356
R779 VAPWR.n69 VAPWR.n67 0.002375
R780 flash_0.x2.clkb flash_0.x2.clkb.t1 167.038
R781 flash_0.x2.clkb flash_0.x2.clkb.t0 87.4292
R782 clk.n1 clk.t2 54.3383
R783 clk.n0 clk.t0 54.3383
R784 clk.n1 clk.t3 53.1307
R785 clk.n0 clk.t1 53.1307
R786 clk.n3 clk 39.2423
R787 clk.n3 clk.n2 9.04175
R788 clk.n2 clk 7.02925
R789 clk.n2 clk 3.72425
R790 clk clk.n1 0.2455
R791 clk clk.n0 0.2455
R792 clk clk.n3 0.078
R793 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t2 649.691
R794 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t0 227.442
R795 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t1 227.361
R796 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t5 216.731
R797 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t6 216.731
R798 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t3 216.731
R799 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t4 216.731
R800 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t7 216.731
R801 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t8 216.731
R802 ui_in[1].n0 ui_in[1].t17 207.43
R803 ui_in[1].n1 ui_in[1].t10 207.43
R804 ui_in[1].n2 ui_in[1].t12 207.43
R805 ui_in[1].n3 ui_in[1].t13 207.43
R806 ui_in[1].n4 ui_in[1].t15 207.43
R807 ui_in[1].n5 ui_in[1].t2 207.43
R808 ui_in[1].n26 ui_in[1].n23 123.867
R809 ui_in[1].n25 ui_in[1] 50.8126
R810 ui_in[1].n15 ui_in[1] 50.8126
R811 ui_in[1] ui_in[1].n1 48.5522
R812 ui_in[1] ui_in[1].n3 48.5522
R813 ui_in[1].n6 ui_in[1].n5 47.7953
R814 ui_in[1].n6 ui_in[1].n2 32.1435
R815 ui_in[1].n8 ui_in[1] 29.9794
R816 ui_in[1].n10 ui_in[1] 29.9794
R817 ui_in[1].n21 ui_in[1] 29.418
R818 ui_in[1].n18 ui_in[1] 29.418
R819 ui_in[1].n27 ui_in[1] 22.2876
R820 ui_in[1].n25 ui_in[1].n24 19.0005
R821 ui_in[1].n21 ui_in[1].n20 19.0005
R822 ui_in[1].n18 ui_in[1].n17 19.0005
R823 ui_in[1].n15 ui_in[1].n14 19.0005
R824 ui_in[1].n8 ui_in[1].n7 19.0005
R825 ui_in[1].n10 ui_in[1].n9 19.0005
R826 ui_in[1] ui_in[1].n0 13.6833
R827 ui_in[1] ui_in[1].n4 13.6833
R828 ui_in[1].n20 ui_in[1].t9 12.0505
R829 ui_in[1].n20 ui_in[1].t6 12.0505
R830 ui_in[1].n17 ui_in[1].t11 12.0505
R831 ui_in[1].n17 ui_in[1].t8 12.0505
R832 ui_in[1].n7 ui_in[1].t5 12.0505
R833 ui_in[1].n7 ui_in[1].t0 12.0505
R834 ui_in[1].n9 ui_in[1].t16 12.0505
R835 ui_in[1].n9 ui_in[1].t14 12.0505
R836 ui_in[1].n27 ui_in[1] 8.72144
R837 ui_in[1].n24 ui_in[1].t3 8.4355
R838 ui_in[1].n24 ui_in[1].t1 8.4355
R839 ui_in[1].n14 ui_in[1].t7 8.4355
R840 ui_in[1].n14 ui_in[1].t4 8.4355
R841 ui_in[1] ui_in[1].n26 4.94473
R842 ui_in[1].n13 ui_in[1].n12 4.5005
R843 ui_in[1].n2 ui_in[1] 3.75222
R844 ui_in[1].n1 ui_in[1] 3.75222
R845 ui_in[1].n0 ui_in[1] 3.75222
R846 ui_in[1].n5 ui_in[1] 3.75222
R847 ui_in[1].n4 ui_in[1] 3.75222
R848 ui_in[1].n3 ui_in[1] 3.75222
R849 ui_in[1].n28 ui_in[1].n13 3.61982
R850 ui_in[1].n11 ui_in[1].n8 2.96269
R851 ui_in[1].n12 ui_in[1].n6 1.69929
R852 ui_in[1].n16 ui_in[1].n15 1.59032
R853 ui_in[1].n22 ui_in[1].n19 1.42722
R854 ui_in[1].n19 ui_in[1].n18 1.32907
R855 ui_in[1].n22 ui_in[1].n21 1.32907
R856 ui_in[1].n26 ui_in[1].n25 1.32907
R857 ui_in[1].n11 ui_in[1].n10 1.32907
R858 ui_in[1].n23 ui_in[1].n16 1.29347
R859 ui_in[1].n12 ui_in[1].n11 0.48697
R860 ui_in[1].n19 ui_in[1].n16 0.25925
R861 ui_in[1].n23 ui_in[1].n22 0.25925
R862 ui_in[1].n13 ui_in[1] 0.0611061
R863 ui_in[1].n28 ui_in[1].n27 0.039875
R864 ui_in[1] ui_in[1].n28 0.0214375
R865 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t2 669.481
R866 flash_0.x4.neg_en_b.n0 flash_0.x4.neg_en_b.t3 669.481
R867 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t0 218.06
R868 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t1 218.06
R869 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t4 211.017
R870 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t6 208.394
R871 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t9 208.394
R872 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t5 207.43
R873 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t7 207.43
R874 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t8 207.43
R875 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.n0 50.3013
R876 flash_0.x4.neg_en_b.n0 flash_0.x4.neg_en_b 29.0914
R877 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t2 649.773
R878 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t3 649.691
R879 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.n1 594.383
R880 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.n2 594.301
R881 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t6 227.361
R882 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t8 216.731
R883 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t14 216.731
R884 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t13 216.731
R885 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t9 105.956
R886 flash_0.x4.neg_mid_b.n0 flash_0.x4.neg_mid_b 103.529
R887 flash_0.x4.neg_mid_b.t8 flash_0.x4.neg_mid_b.t7 101.221
R888 flash_0.x4.neg_mid_b.t14 flash_0.x4.neg_mid_b.t12 101.221
R889 flash_0.x4.neg_mid_b.t13 flash_0.x4.neg_mid_b.t11 101.221
R890 flash_0.x4.neg_mid_b.n1 flash_0.x4.neg_mid_b.t4 55.3905
R891 flash_0.x4.neg_mid_b.n1 flash_0.x4.neg_mid_b.t5 55.3905
R892 flash_0.x4.neg_mid_b.n2 flash_0.x4.neg_mid_b.t1 55.3905
R893 flash_0.x4.neg_mid_b.n2 flash_0.x4.neg_mid_b.t0 55.3905
R894 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.n0 23.6062
R895 flash_0.x4.neg_mid_b.n0 flash_0.x4.neg_mid_b.t10 22.3887
R896 flash_0.x4.VOUT flash_0.x4.VOUT.t4 649.691
R897 flash_0.x4.VOUT flash_0.x4.VOUT.t1 649.691
R898 flash_0.x4.VOUT flash_0.x4.VOUT.t12 649.691
R899 flash_0.x4.VOUT flash_0.x4.VOUT.t8 649.691
R900 flash_0.x4.VOUT flash_0.x4.VOUT.n0 594.383
R901 flash_0.x4.VOUT flash_0.x4.VOUT.n3 594.301
R902 flash_0.x4.VOUT flash_0.x4.VOUT.n1 594.301
R903 flash_0.x4.VOUT flash_0.x4.VOUT.n2 594.301
R904 flash_0.x4.VOUT flash_0.x4.VOUT.t7 227.431
R905 flash_0.x4.VOUT flash_0.x4.VOUT.t0 227.361
R906 flash_0.x4.VOUT flash_0.x4.VOUT.t14 149.423
R907 flash_0.x4.VOUT.n3 flash_0.x4.VOUT.t2 55.3905
R908 flash_0.x4.VOUT.n3 flash_0.x4.VOUT.t5 55.3905
R909 flash_0.x4.VOUT.n1 flash_0.x4.VOUT.t13 55.3905
R910 flash_0.x4.VOUT.n1 flash_0.x4.VOUT.t9 55.3905
R911 flash_0.x4.VOUT.n0 flash_0.x4.VOUT.t11 55.3905
R912 flash_0.x4.VOUT.n0 flash_0.x4.VOUT.t10 55.3905
R913 flash_0.x4.VOUT.n2 flash_0.x4.VOUT.t6 55.3905
R914 flash_0.x4.VOUT.n2 flash_0.x4.VOUT.t3 55.3905
R915 flash_0.x4.dcgint.n0 flash_0.x4.dcgint.t5 644.461
R916 flash_0.x4.dcgint.n5 flash_0.x4.dcgint.t3 640.39
R917 flash_0.x4.dcgint.n3 flash_0.x4.dcgint.n1 605.365
R918 flash_0.x4.dcgint.n3 flash_0.x4.dcgint.n2 605.365
R919 flash_0.x4.dcgint.n4 flash_0.x4.dcgint.t2 477.228
R920 flash_0.x4.dcgint.t2 flash_0.x4.dcgint.t0 339.594
R921 flash_0.x4.dcgint.t0 flash_0.x4.dcgint.t6 339.594
R922 flash_0.x4.dcgint flash_0.x4.dcgint.t11 227.361
R923 flash_0.x4.dcgint flash_0.x4.dcgint.t10 227.361
R924 flash_0.x4.dcgint flash_0.x4.dcgint.t9 227.361
R925 flash_0.x4.dcgint.n4 flash_0.x4.dcgint.n3 69.5657
R926 flash_0.x4.dcgint.n1 flash_0.x4.dcgint.t1 55.3905
R927 flash_0.x4.dcgint.n1 flash_0.x4.dcgint.t7 55.3905
R928 flash_0.x4.dcgint.n2 flash_0.x4.dcgint.t4 55.3905
R929 flash_0.x4.dcgint.n2 flash_0.x4.dcgint.t8 55.3905
R930 flash_0.x4.dcgint.n6 flash_0.x4.dcgint.n5 9.3005
R931 flash_0.x4.dcgint.n5 flash_0.x4.dcgint.n4 8.9605
R932 flash_0.x4.dcgint flash_0.x4.dcgint.n6 7.52362
R933 flash_0.x4.dcgint.n6 flash_0.x4.dcgint.n0 1.14684
R934 flash_0.x4.dcgint.n4 flash_0.x4.dcgint.n0 1.0086
R935 flash_0.x7.pos_en_b.n1 flash_0.x7.pos_en_b.t3 669.481
R936 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b.t0 669.481
R937 flash_0.x7.pos_en_b flash_0.x7.pos_en_b.t1 218.06
R938 flash_0.x7.pos_en_b flash_0.x7.pos_en_b.t2 218.06
R939 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b.t6 65.4032
R940 flash_0.x7.pos_en_b.t6 flash_0.x7.pos_en_b 56.2429
R941 flash_0.x7.pos_en_b.t6 flash_0.x7.pos_en_b 56.2429
R942 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b 50.8126
R943 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b 50.8126
R944 flash_0.x7.pos_en_b flash_0.x7.pos_en_b.n1 29.0914
R945 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b 29.0914
R946 flash_0.x7.pos_en_b.n1 flash_0.x7.pos_en_b.n0 28.2591
R947 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b.t4 27.4355
R948 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b.t5 27.4355
R949 VDPWR.n84 VDPWR.n70 5586
R950 VDPWR.n84 VDPWR.n71 5586
R951 VDPWR.n79 VDPWR.n71 5586
R952 VDPWR.n79 VDPWR.n70 5586
R953 VDPWR.n129 VDPWR.n115 5586
R954 VDPWR.n129 VDPWR.n116 5586
R955 VDPWR.n124 VDPWR.n116 5586
R956 VDPWR.n124 VDPWR.n115 5586
R957 VDPWR.n30 VDPWR.n29 4689.72
R958 VDPWR.n27 VDPWR.n25 4689.72
R959 VDPWR.n80 VDPWR.n72 4509.29
R960 VDPWR.n125 VDPWR.n117 4509.29
R961 VDPWR.n83 VDPWR.n72 4506
R962 VDPWR.n128 VDPWR.n117 4506
R963 VDPWR.n44 VDPWR.n37 2442.35
R964 VDPWR.n41 VDPWR.n38 2442.35
R965 VDPWR.n61 VDPWR.n54 2442.35
R966 VDPWR.n58 VDPWR.n55 2442.35
R967 VDPWR.n83 VDPWR.t29 2271.78
R968 VDPWR.n128 VDPWR.t37 2271.78
R969 VDPWR.n30 VDPWR.n24 1828.1
R970 VDPWR.n28 VDPWR.n27 1828.1
R971 VDPWR.t0 VDPWR.t42 1429.17
R972 VDPWR.t40 VDPWR.t25 1429.17
R973 VDPWR.t29 VDPWR.n82 1226.56
R974 VDPWR.t37 VDPWR.n127 1226.56
R975 VDPWR.n26 VDPWR.n22 902.777
R976 VDPWR.n26 VDPWR.n23 902.777
R977 VDPWR.n31 VDPWR.n23 881.453
R978 VDPWR.n32 VDPWR.n22 879.466
R979 VDPWR.n33 VDPWR.t46 649.831
R980 VDPWR.n85 VDPWR.n69 627.201
R981 VDPWR.n78 VDPWR.n68 627.201
R982 VDPWR.n130 VDPWR.n114 627.201
R983 VDPWR.n123 VDPWR.n113 627.201
R984 VDPWR.n103 VDPWR.n102 585
R985 VDPWR.n98 VDPWR.n97 585
R986 VDPWR.n93 VDPWR.n92 585
R987 VDPWR.n101 VDPWR.n100 585
R988 VDPWR.n96 VDPWR.n95 585
R989 VDPWR.n91 VDPWR.n90 585
R990 VDPWR.n14 VDPWR.n13 585
R991 VDPWR.n9 VDPWR.n8 585
R992 VDPWR.n4 VDPWR.n3 585
R993 VDPWR.n12 VDPWR.n11 585
R994 VDPWR.n7 VDPWR.n6 585
R995 VDPWR.n2 VDPWR.n1 585
R996 VDPWR.n42 VDPWR.n37 535.419
R997 VDPWR.n43 VDPWR.n38 535.419
R998 VDPWR.n59 VDPWR.n54 535.419
R999 VDPWR.n60 VDPWR.n55 535.419
R1000 VDPWR.n86 VDPWR.n85 525.553
R1001 VDPWR.n131 VDPWR.n130 525.553
R1002 VDPWR.n77 VDPWR.n69 492.048
R1003 VDPWR.n122 VDPWR.n114 492.048
R1004 VDPWR.n82 VDPWR.t0 394.779
R1005 VDPWR.n127 VDPWR.t40 394.779
R1006 VDPWR.n88 VDPWR.n66 297.151
R1007 VDPWR.n107 VDPWR.n106 297.151
R1008 VDPWR.n18 VDPWR.n17 297.151
R1009 VDPWR.n111 VDPWR.n0 297.151
R1010 VDPWR.n81 VDPWR.t20 272.363
R1011 VDPWR.n126 VDPWR.t47 272.363
R1012 VDPWR.n40 VDPWR.n36 260.519
R1013 VDPWR.n45 VDPWR.n36 260.519
R1014 VDPWR.n57 VDPWR.n53 260.519
R1015 VDPWR.n62 VDPWR.n53 260.519
R1016 VDPWR.n40 VDPWR.n39 232.66
R1017 VDPWR.n46 VDPWR.n45 232.66
R1018 VDPWR.n57 VDPWR.n56 232.66
R1019 VDPWR.n63 VDPWR.n62 232.66
R1020 VDPWR.n34 VDPWR.t54 228.215
R1021 VDPWR.n51 VDPWR.t5 228.215
R1022 VDPWR.t14 VDPWR.t22 172.133
R1023 VDPWR.t12 VDPWR.t16 172.133
R1024 VDPWR.t18 VDPWR.t12 172.133
R1025 VDPWR.t20 VDPWR.t18 172.133
R1026 VDPWR.t27 VDPWR.t6 172.133
R1027 VDPWR.t51 VDPWR.t2 172.133
R1028 VDPWR.t9 VDPWR.t51 172.133
R1029 VDPWR.t47 VDPWR.t9 172.133
R1030 VDPWR.n66 VDPWR.t1 160.44
R1031 VDPWR.n66 VDPWR.t30 160.44
R1032 VDPWR.n106 VDPWR.t33 160.44
R1033 VDPWR.n106 VDPWR.t43 160.44
R1034 VDPWR.n17 VDPWR.t50 160.44
R1035 VDPWR.n17 VDPWR.t26 160.44
R1036 VDPWR.n0 VDPWR.t41 160.44
R1037 VDPWR.n0 VDPWR.t38 160.44
R1038 VDPWR.n78 VDPWR.n77 135.154
R1039 VDPWR.n123 VDPWR.n122 135.154
R1040 VDPWR.t32 VDPWR.t14 135.093
R1041 VDPWR.t49 VDPWR.t27 135.093
R1042 VDPWR.n74 VDPWR 106.918
R1043 VDPWR.n119 VDPWR 106.918
R1044 VDPWR.n86 VDPWR.n68 101.647
R1045 VDPWR.n131 VDPWR.n113 101.647
R1046 VDPWR.n81 VDPWR.n80 57.7708
R1047 VDPWR.n126 VDPWR.n125 57.7708
R1048 VDPWR.n102 VDPWR.t31 55.3905
R1049 VDPWR.n102 VDPWR.t21 55.3905
R1050 VDPWR.n97 VDPWR.t17 55.3905
R1051 VDPWR.n97 VDPWR.t39 55.3905
R1052 VDPWR.n92 VDPWR.t36 55.3905
R1053 VDPWR.n92 VDPWR.t15 55.3905
R1054 VDPWR.n100 VDPWR.t19 55.3905
R1055 VDPWR.n100 VDPWR.t35 55.3905
R1056 VDPWR.n95 VDPWR.t34 55.3905
R1057 VDPWR.n95 VDPWR.t13 55.3905
R1058 VDPWR.n90 VDPWR.t23 55.3905
R1059 VDPWR.n90 VDPWR.t44 55.3905
R1060 VDPWR.n13 VDPWR.t10 55.3905
R1061 VDPWR.n13 VDPWR.t48 55.3905
R1062 VDPWR.n8 VDPWR.t8 55.3905
R1063 VDPWR.n8 VDPWR.t55 55.3905
R1064 VDPWR.n3 VDPWR.t11 55.3905
R1065 VDPWR.n3 VDPWR.t28 55.3905
R1066 VDPWR.n11 VDPWR.t24 55.3905
R1067 VDPWR.n11 VDPWR.t57 55.3905
R1068 VDPWR.n6 VDPWR.t3 55.3905
R1069 VDPWR.n6 VDPWR.t52 55.3905
R1070 VDPWR.n1 VDPWR.t7 55.3905
R1071 VDPWR.n1 VDPWR.t56 55.3905
R1072 VDPWR.t16 VDPWR.t32 37.0418
R1073 VDPWR.t2 VDPWR.t49 37.0418
R1074 VDPWR.n27 VDPWR.n26 37.0005
R1075 VDPWR.n31 VDPWR.n30 37.0005
R1076 VDPWR.n38 VDPWR.n36 30.8338
R1077 VDPWR.n37 VDPWR.n35 30.8338
R1078 VDPWR.n55 VDPWR.n53 30.8338
R1079 VDPWR.n54 VDPWR.n52 30.8338
R1080 VDPWR.n39 VDPWR.n35 27.8593
R1081 VDPWR.n46 VDPWR.n35 27.8593
R1082 VDPWR.n56 VDPWR.n52 27.8593
R1083 VDPWR.n63 VDPWR.n52 27.8593
R1084 VDPWR.n74 VDPWR.n73 19.0005
R1085 VDPWR.n119 VDPWR.n118 19.0005
R1086 VDPWR.n41 VDPWR.n40 16.8187
R1087 VDPWR.n45 VDPWR.n44 16.8187
R1088 VDPWR.n58 VDPWR.n57 16.8187
R1089 VDPWR.n62 VDPWR.n61 16.8187
R1090 VDPWR.n103 VDPWR 14.3064
R1091 VDPWR.n98 VDPWR 14.3064
R1092 VDPWR.n93 VDPWR 14.3064
R1093 VDPWR.n101 VDPWR 14.3064
R1094 VDPWR.n96 VDPWR 14.3064
R1095 VDPWR.n91 VDPWR 14.3064
R1096 VDPWR.n14 VDPWR 14.3064
R1097 VDPWR.n9 VDPWR 14.3064
R1098 VDPWR.n4 VDPWR 14.3064
R1099 VDPWR.n12 VDPWR 14.3064
R1100 VDPWR.n7 VDPWR 14.3064
R1101 VDPWR.n2 VDPWR 14.3064
R1102 VDPWR.n104 VDPWR.n103 13.8019
R1103 VDPWR.n99 VDPWR.n98 13.8019
R1104 VDPWR.n94 VDPWR.n93 13.8019
R1105 VDPWR.n104 VDPWR.n101 13.8019
R1106 VDPWR.n99 VDPWR.n96 13.8019
R1107 VDPWR.n94 VDPWR.n91 13.8019
R1108 VDPWR.n15 VDPWR.n14 13.8019
R1109 VDPWR.n10 VDPWR.n9 13.8019
R1110 VDPWR.n5 VDPWR.n4 13.8019
R1111 VDPWR.n15 VDPWR.n12 13.8019
R1112 VDPWR.n10 VDPWR.n7 13.8019
R1113 VDPWR.n5 VDPWR.n2 13.8019
R1114 VDPWR.n42 VDPWR.n41 13.0425
R1115 VDPWR.n44 VDPWR.n43 13.0425
R1116 VDPWR.n59 VDPWR.n58 13.0425
R1117 VDPWR.n61 VDPWR.n60 13.0425
R1118 VDPWR.t42 VDPWR.n81 10.895
R1119 VDPWR.t25 VDPWR.n126 10.895
R1120 VDPWR.n85 VDPWR.n84 10.2783
R1121 VDPWR.n84 VDPWR.n83 10.2783
R1122 VDPWR.n79 VDPWR.n78 10.2783
R1123 VDPWR.n80 VDPWR.n79 10.2783
R1124 VDPWR.n130 VDPWR.n129 10.2783
R1125 VDPWR.n129 VDPWR.n128 10.2783
R1126 VDPWR.n124 VDPWR.n123 10.2783
R1127 VDPWR.n125 VDPWR.n124 10.2783
R1128 VDPWR.n65 VDPWR.n64 9.74376
R1129 VDPWR.n39 VDPWR.n34 9.35589
R1130 VDPWR.n56 VDPWR.n51 9.35589
R1131 VDPWR VDPWR.n46 9.33194
R1132 VDPWR VDPWR.n63 9.33194
R1133 VDPWR.n73 VDPWR.t59 8.4355
R1134 VDPWR.n73 VDPWR.t58 8.4355
R1135 VDPWR.n118 VDPWR.t61 8.4355
R1136 VDPWR.n118 VDPWR.t60 8.4355
R1137 VDPWR.n70 VDPWR.n69 6.37981
R1138 VDPWR.n72 VDPWR.n70 6.37981
R1139 VDPWR.n71 VDPWR.n68 6.37981
R1140 VDPWR.n82 VDPWR.n71 6.37981
R1141 VDPWR.n115 VDPWR.n114 6.37981
R1142 VDPWR.n117 VDPWR.n115 6.37981
R1143 VDPWR.n116 VDPWR.n113 6.37981
R1144 VDPWR.n127 VDPWR.n116 6.37981
R1145 VDPWR.n48 VDPWR.n33 5.59737
R1146 VDPWR.n75 VDPWR.n67 4.51137
R1147 VDPWR.n120 VDPWR.n112 4.51137
R1148 VDPWR.n111 VDPWR.n110 3.96097
R1149 VDPWR.n89 VDPWR.n88 3.9605
R1150 VDPWR.n77 VDPWR.n76 3.88885
R1151 VDPWR.n122 VDPWR.n121 3.88885
R1152 VDPWR.n20 VDPWR 3.84311
R1153 VDPWR.n87 VDPWR.n67 3.7551
R1154 VDPWR.n132 VDPWR.n112 3.7551
R1155 VDPWR.n43 VDPWR.t53 3.68792
R1156 VDPWR.t53 VDPWR.n42 3.68792
R1157 VDPWR.n60 VDPWR.t4 3.68792
R1158 VDPWR.t4 VDPWR.n59 3.68792
R1159 VDPWR.n25 VDPWR.n22 3.03329
R1160 VDPWR.n29 VDPWR.n23 3.03329
R1161 VDPWR.n76 VDPWR.n74 2.3749
R1162 VDPWR.n121 VDPWR.n119 2.3749
R1163 VDPWR.n19 VDPWR.n18 2.25658
R1164 VDPWR.n108 VDPWR.n107 2.2555
R1165 VDPWR.n110 VDPWR.n19 1.98603
R1166 VDPWR.n33 VDPWR.n32 1.8605
R1167 VDPWR.n25 VDPWR.n24 1.85038
R1168 VDPWR.n29 VDPWR.n28 1.85038
R1169 VDPWR.n109 VDPWR.n108 1.7055
R1170 VDPWR.n49 VDPWR.n48 1.43592
R1171 VDPWR.n65 VDPWR.n50 1.29333
R1172 VDPWR.n28 VDPWR.t45 1.18321
R1173 VDPWR.t45 VDPWR.n24 1.18321
R1174 VDPWR.n32 VDPWR.n31 1.0245
R1175 VDPWR.n76 VDPWR.n75 0.813
R1176 VDPWR.n121 VDPWR.n120 0.813
R1177 VDPWR.n89 VDPWR.n65 0.683034
R1178 VDPWR.n85 VDPWR.n67 0.547559
R1179 VDPWR.n130 VDPWR.n112 0.547559
R1180 VDPWR.n48 VDPWR.n47 0.53175
R1181 VDPWR.n50 VDPWR.n49 0.486785
R1182 VDPWR.n110 VDPWR.n109 0.475641
R1183 VDPWR.n87 VDPWR.n86 0.4655
R1184 VDPWR.n132 VDPWR.n131 0.4655
R1185 VDPWR.n75 VDPWR.n69 0.344944
R1186 VDPWR.n120 VDPWR.n114 0.344944
R1187 VDPWR.n109 VDPWR.n89 0.278606
R1188 VDPWR.n19 VDPWR.n16 0.201021
R1189 VDPWR.n108 VDPWR.n105 0.182167
R1190 VDPWR.n21 VDPWR.n20 0.171
R1191 VDPWR.n107 VDPWR 0.102773
R1192 VDPWR.n18 VDPWR 0.102773
R1193 VDPWR.n99 VDPWR.n94 0.0902727
R1194 VDPWR.n10 VDPWR.n5 0.0902727
R1195 VDPWR.n105 VDPWR.n99 0.0772045
R1196 VDPWR.n16 VDPWR.n10 0.0772045
R1197 VDPWR.n21 VDPWR 0.0558125
R1198 VDPWR.n50 VDPWR.n20 0.0483835
R1199 VDPWR.n88 VDPWR 0.0483723
R1200 VDPWR VDPWR.n111 0.0483723
R1201 VDPWR.n47 VDPWR 0.0199611
R1202 VDPWR.n64 VDPWR 0.0199611
R1203 VDPWR.n49 VDPWR.n21 0.014875
R1204 VDPWR.n105 VDPWR.n104 0.0135682
R1205 VDPWR.n16 VDPWR.n15 0.0135682
R1206 VDPWR.n47 VDPWR.n34 0.00499102
R1207 VDPWR.n64 VDPWR.n51 0.00499102
R1208 VDPWR VDPWR.n87 0.00116489
R1209 VDPWR VDPWR.n132 0.00116489
R1210 ua[0].n6 ua[0].n4 2724.21
R1211 ua[0].n9 ua[0].n8 2724.21
R1212 ua[0].n7 ua[0].n6 1018.07
R1213 ua[0].n9 ua[0].n3 1018.07
R1214 ua[0].n12 ua[0].t1 649.886
R1215 ua[0].n0 ua[0].t3 649.692
R1216 ua[0].n5 ua[0].n1 526.307
R1217 ua[0].n5 ua[0].n2 526.307
R1218 ua[0].n10 ua[0].n2 497.486
R1219 ua[0].n11 ua[0].n1 493.762
R1220 ua[0].n6 ua[0].n5 37.0005
R1221 ua[0].n10 ua[0].n9 37.0005
R1222 ua[0].n14 ua[0] 13.435
R1223 ua[0].n4 ua[0].n1 5.78175
R1224 ua[0].n8 ua[0].n2 5.78175
R1225 ua[0].n0 ua[0].t2 4.69622
R1226 ua[0].n4 ua[0].n3 3.61407
R1227 ua[0].n8 ua[0].n7 3.61407
R1228 ua[0].t0 ua[0].n3 2.16152
R1229 ua[0].n7 ua[0].t0 2.16152
R1230 ua[0].n12 ua[0].n11 1.8605
R1231 ua[0].n11 ua[0].n10 1.54533
R1232 ua[0].n14 ua[0].n13 0.9005
R1233 ua[0].n13 ua[0].n0 0.64055
R1234 ua[0].n13 ua[0].n12 0.405262
R1235 ua[0] ua[0].n14 0.0639375
R1236 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t2 669.481
R1237 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t1 669.481
R1238 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t3 218.06
R1239 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t0 218.06
R1240 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t9 211.017
R1241 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t8 208.394
R1242 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t6 208.394
R1243 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t4 207.43
R1244 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t7 207.43
R1245 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t5 207.43
R1246 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t0 649.773
R1247 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t5 649.691
R1248 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.n3 594.383
R1249 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.n4 594.301
R1250 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t6 227.361
R1251 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t8 216.731
R1252 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t13 216.731
R1253 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t14 216.731
R1254 flash_0.x7.neg_mid_b.n0 flash_0.x7.neg_mid_b.t15 105.956
R1255 flash_0.x7.neg_mid_b.n2 flash_0.x7.neg_mid_b 103.529
R1256 flash_0.x7.neg_mid_b.t8 flash_0.x7.neg_mid_b.t7 101.221
R1257 flash_0.x7.neg_mid_b.t13 flash_0.x7.neg_mid_b.t11 101.221
R1258 flash_0.x7.neg_mid_b.t14 flash_0.x7.neg_mid_b.t12 101.221
R1259 flash_0.x7.neg_mid_b.n4 flash_0.x7.neg_mid_b.t4 55.3905
R1260 flash_0.x7.neg_mid_b.n4 flash_0.x7.neg_mid_b.t2 55.3905
R1261 flash_0.x7.neg_mid_b.n3 flash_0.x7.neg_mid_b.t3 55.3905
R1262 flash_0.x7.neg_mid_b.n3 flash_0.x7.neg_mid_b.t1 55.3905
R1263 flash_0.x7.neg_mid_b.n2 flash_0.x7.neg_mid_b.n1 22.3887
R1264 flash_0.x7.neg_mid_b.n1 flash_0.x7.neg_mid_b.t10 8.4355
R1265 flash_0.x7.neg_mid_b.n1 flash_0.x7.neg_mid_b.t9 8.4355
R1266 flash_0.x7.neg_mid_b.n0 flash_0.x7.neg_mid_b 5.14452
R1267 flash_0.x7.neg_mid_b.n0 flash_0.x7.neg_mid_b.n2 2.45104
R1268 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.n0 1.98963
R1269 flash_0.x6.Y flash_0.x6.Y.t0 84.4155
R1270 flash_0.x5.A.n6 flash_0.x5.A.n4 2888.05
R1271 flash_0.x5.A.n9 flash_0.x5.A.n3 2888.05
R1272 flash_0.x5.A.n11 flash_0.x5.A.t0 658.039
R1273 flash_0.x5.A.n8 flash_0.x5.A.n4 509.978
R1274 flash_0.x5.A.n7 flash_0.x5.A.n3 509.978
R1275 flash_0.x5.A.n5 flash_0.x5.A.n2 334.683
R1276 flash_0.x5.A.n10 flash_0.x5.A.n2 334.683
R1277 flash_0.x5.A.n5 flash_0.x5.A.n1 291.084
R1278 flash_0.x5.A.n1 flash_0.x5.A.n10 290.635
R1279 flash_0.x5.A.n0 flash_0.x5.A.t1 215.056
R1280 flash_0.x5.A.n6 flash_0.x5.A.n5 146.25
R1281 flash_0.x5.A.n10 flash_0.x5.A.n9 146.25
R1282 flash_0.x5.A.n7 flash_0.x5.A.n6 114.621
R1283 flash_0.x5.A.n9 flash_0.x5.A.n8 114.621
R1284 flash_0.x5.A flash_0.x5.A.t4 33.6612
R1285 flash_0.x5.A flash_0.x5.A.t5 32.9049
R1286 flash_0.x5.A.n4 flash_0.x5.A.n2 32.5005
R1287 flash_0.x5.A.n3 flash_0.x5.A.n1 32.5005
R1288 flash_0.x5.A.t2 flash_0.x5.A.n7 25.8261
R1289 flash_0.x5.A.n8 flash_0.x5.A.t2 25.8261
R1290 flash_0.x5.A.n0 flash_0.x5.A.t3 17.2847
R1291 flash_0.x5.A flash_0.x5.A.n11 2.49814
R1292 flash_0.x5.A.n0 flash_0.x5.A.n1 1.43573
R1293 flash_0.x5.A.n11 flash_0.x5.A.n0 1.12981
R1294 ui_in[0].n0 ui_in[0].t6 207.43
R1295 ui_in[0].n1 ui_in[0].t14 207.43
R1296 ui_in[0].n2 ui_in[0].t8 207.43
R1297 ui_in[0].n3 ui_in[0].t9 207.43
R1298 ui_in[0].n4 ui_in[0].t0 207.43
R1299 ui_in[0].n5 ui_in[0].t10 207.43
R1300 ui_in[0].n26 ui_in[0].n23 123.867
R1301 ui_in[0].n25 ui_in[0] 50.8126
R1302 ui_in[0].n15 ui_in[0] 50.8126
R1303 ui_in[0] ui_in[0].n1 48.5522
R1304 ui_in[0] ui_in[0].n3 48.5522
R1305 ui_in[0].n6 ui_in[0].n5 47.7953
R1306 ui_in[0].n6 ui_in[0].n2 32.1435
R1307 ui_in[0].n8 ui_in[0] 29.9794
R1308 ui_in[0].n10 ui_in[0] 29.9794
R1309 ui_in[0].n21 ui_in[0] 29.418
R1310 ui_in[0].n18 ui_in[0] 29.418
R1311 ui_in[0].n27 ui_in[0] 26.7297
R1312 ui_in[0].n25 ui_in[0].n24 19.0005
R1313 ui_in[0].n21 ui_in[0].n20 19.0005
R1314 ui_in[0].n18 ui_in[0].n17 19.0005
R1315 ui_in[0].n15 ui_in[0].n14 19.0005
R1316 ui_in[0].n8 ui_in[0].n7 19.0005
R1317 ui_in[0].n10 ui_in[0].n9 19.0005
R1318 ui_in[0] ui_in[0].n0 13.6833
R1319 ui_in[0] ui_in[0].n4 13.6833
R1320 ui_in[0].n20 ui_in[0].t17 12.0505
R1321 ui_in[0].n20 ui_in[0].t15 12.0505
R1322 ui_in[0].n17 ui_in[0].t7 12.0505
R1323 ui_in[0].n17 ui_in[0].t4 12.0505
R1324 ui_in[0].n7 ui_in[0].t16 12.0505
R1325 ui_in[0].n7 ui_in[0].t12 12.0505
R1326 ui_in[0].n9 ui_in[0].t5 12.0505
R1327 ui_in[0].n9 ui_in[0].t2 12.0505
R1328 ui_in[0] ui_in[0].n13 11.4683
R1329 ui_in[0].n24 ui_in[0].t13 8.4355
R1330 ui_in[0].n24 ui_in[0].t11 8.4355
R1331 ui_in[0].n14 ui_in[0].t3 8.4355
R1332 ui_in[0].n14 ui_in[0].t1 8.4355
R1333 ui_in[0] ui_in[0].n26 4.94473
R1334 ui_in[0].n13 ui_in[0].n12 4.5005
R1335 ui_in[0].n13 ui_in[0] 4.0005
R1336 ui_in[0].n2 ui_in[0] 3.75222
R1337 ui_in[0].n1 ui_in[0] 3.75222
R1338 ui_in[0].n0 ui_in[0] 3.75222
R1339 ui_in[0].n5 ui_in[0] 3.75222
R1340 ui_in[0].n4 ui_in[0] 3.75222
R1341 ui_in[0].n3 ui_in[0] 3.75222
R1342 ui_in[0].n11 ui_in[0].n8 2.96269
R1343 ui_in[0].n27 ui_in[0] 2.12895
R1344 ui_in[0].n12 ui_in[0].n6 1.69929
R1345 ui_in[0].n16 ui_in[0].n15 1.59032
R1346 ui_in[0].n22 ui_in[0].n19 1.42722
R1347 ui_in[0].n19 ui_in[0].n18 1.32907
R1348 ui_in[0].n22 ui_in[0].n21 1.32907
R1349 ui_in[0].n26 ui_in[0].n25 1.32907
R1350 ui_in[0].n11 ui_in[0].n10 1.32907
R1351 ui_in[0].n23 ui_in[0].n16 1.29347
R1352 ui_in[0].n12 ui_in[0].n11 0.48697
R1353 ui_in[0].n19 ui_in[0].n16 0.25925
R1354 ui_in[0].n23 ui_in[0].n22 0.25925
R1355 ui_in[0].n13 ui_in[0] 0.0611061
R1356 ui_in[0] ui_in[0].n27 0.02925
R1357 flash_0.x7.VOUT.n8 flash_0.x7.VOUT.n6 2045.32
R1358 flash_0.x7.VOUT.n11 flash_0.x7.VOUT.n5 2045.32
R1359 flash_0.x7.VOUT.n9 flash_0.x7.VOUT.n8 836.909
R1360 flash_0.x7.VOUT.n11 flash_0.x7.VOUT.n10 836.909
R1361 flash_0.x7.VOUT flash_0.x7.VOUT.t5 649.691
R1362 flash_0.x7.VOUT flash_0.x7.VOUT.t12 649.691
R1363 flash_0.x7.VOUT flash_0.x7.VOUT.t11 649.691
R1364 flash_0.x7.VOUT flash_0.x7.VOUT.t7 649.691
R1365 flash_0.x7.VOUT flash_0.x7.VOUT.n2 594.383
R1366 flash_0.x7.VOUT flash_0.x7.VOUT.n13 594.301
R1367 flash_0.x7.VOUT flash_0.x7.VOUT.n14 594.301
R1368 flash_0.x7.VOUT flash_0.x7.VOUT.n3 594.301
R1369 flash_0.x7.VOUT flash_0.x7.VOUT.t0 227.431
R1370 flash_0.x7.VOUT flash_0.x7.VOUT.t1 227.361
R1371 flash_0.x7.VOUT.n6 flash_0.x7.VOUT.n4 195
R1372 flash_0.x7.VOUT.n12 flash_0.x7.VOUT.n11 146.25
R1373 flash_0.x7.VOUT.n8 flash_0.x7.VOUT.n7 146.25
R1374 flash_0.x7.VOUT.n12 flash_0.x7.VOUT.n4 132.894
R1375 flash_0.x7.VOUT.n7 flash_0.x7.VOUT.n4 132.894
R1376 flash_0.x7.VOUT.n9 flash_0.x7.VOUT.n5 105.183
R1377 flash_0.x7.VOUT.n10 flash_0.x7.VOUT.n6 105.183
R1378 flash_0.x7.VOUT.n12 flash_0.x7.VOUT.n1 53.1377
R1379 flash_0.x7.VOUT.n10 flash_0.x7.VOUT.t14 79.7913
R1380 flash_0.x7.VOUT.t14 flash_0.x7.VOUT.n9 79.7913
R1381 flash_0.x7.VOUT.n13 flash_0.x7.VOUT.t6 55.3905
R1382 flash_0.x7.VOUT.n13 flash_0.x7.VOUT.t4 55.3905
R1383 flash_0.x7.VOUT.n14 flash_0.x7.VOUT.t2 55.3905
R1384 flash_0.x7.VOUT.n14 flash_0.x7.VOUT.t3 55.3905
R1385 flash_0.x7.VOUT.n3 flash_0.x7.VOUT.t8 55.3905
R1386 flash_0.x7.VOUT.n3 flash_0.x7.VOUT.t9 55.3905
R1387 flash_0.x7.VOUT.n2 flash_0.x7.VOUT.t13 55.3905
R1388 flash_0.x7.VOUT.n2 flash_0.x7.VOUT.t10 55.3905
R1389 flash_0.x7.VOUT.n7 flash_0.x7.VOUT.n0 52.7987
R1390 flash_0.x7.VOUT flash_0.x7.VOUT.n0 28.5614
R1391 flash_0.x7.VOUT.n0 flash_0.x7.VOUT.n1 0.446827
R1392 flash_0.x7.VOUT.n5 flash_0.x7.VOUT.n1 198.951
R1393 w_7728_24730.t0 w_7728_24730.t2 336.07
R1394 w_7728_24730.t3 w_7728_24730.t0 649.856
R1395 w_7728_24730.t0 w_7728_24730.t1 649.692
R1396 flash_0.x3.clka flash_0.x3.clka.t1 167.038
R1397 flash_0.x3.clka flash_0.x3.clka.t0 87.4292
R1398 flash_0.x3.clkb flash_0.x3.clkb.t1 167.038
R1399 flash_0.x3.clkb flash_0.x3.clkb.t0 87.4292
R1400 flash_0.x4.pos_en_b.n0 flash_0.x4.pos_en_b.t0 669.481
R1401 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.t1 669.481
R1402 flash_0.x4.pos_en_b flash_0.x4.pos_en_b.t3 218.06
R1403 flash_0.x4.pos_en_b flash_0.x4.pos_en_b.t2 218.06
R1404 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.t4 65.4032
R1405 flash_0.x4.pos_en_b.t4 flash_0.x4.pos_en_b 56.2429
R1406 flash_0.x4.pos_en_b.t4 flash_0.x4.pos_en_b 56.2429
R1407 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b 50.8126
R1408 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b 50.8126
R1409 flash_0.x4.pos_en_b flash_0.x4.pos_en_b.n1 29.0914
R1410 flash_0.x4.pos_en_b.n0 flash_0.x4.pos_en_b 29.0914
R1411 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.n0 28.2591
R1412 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.t5 27.4355
R1413 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.t6 27.4355
R1414 ui_in[2].n1 ui_in[2].t1 150.088
R1415 ui_in[2].n0 ui_in[2].t2 33.6007
R1416 ui_in[2].n0 ui_in[2].t0 32.9049
R1417 ui_in[2].n2 ui_in[2] 31.3871
R1418 ui_in[2].n2 ui_in[2].n1 4.55612
R1419 ui_in[2].n1 ui_in[2] 1.9712
R1420 ui_in[2] ui_in[2].n0 0.063
R1421 ui_in[2] ui_in[2].n2 0.047375
R1422 flash_0.x2.clka flash_0.x2.clka.t1 167.038
R1423 flash_0.x2.clka flash_0.x2.clka.t0 87.4292
R1424 flash_0.x7.dcgint.n0 flash_0.x7.dcgint.t7 644.461
R1425 flash_0.x7.dcgint.n5 flash_0.x7.dcgint.t4 640.39
R1426 flash_0.x7.dcgint.n3 flash_0.x7.dcgint.n1 605.365
R1427 flash_0.x7.dcgint.n3 flash_0.x7.dcgint.n2 605.365
R1428 flash_0.x7.dcgint.n4 flash_0.x7.dcgint.t3 477.228
R1429 flash_0.x7.dcgint.t3 flash_0.x7.dcgint.t5 339.594
R1430 flash_0.x7.dcgint.t5 flash_0.x7.dcgint.t9 339.594
R1431 flash_0.x7.dcgint flash_0.x7.dcgint.t2 227.361
R1432 flash_0.x7.dcgint flash_0.x7.dcgint.t1 227.361
R1433 flash_0.x7.dcgint flash_0.x7.dcgint.t0 227.361
R1434 flash_0.x7.dcgint.n4 flash_0.x7.dcgint.n3 69.5657
R1435 flash_0.x7.dcgint.n1 flash_0.x7.dcgint.t6 55.3905
R1436 flash_0.x7.dcgint.n1 flash_0.x7.dcgint.t10 55.3905
R1437 flash_0.x7.dcgint.n2 flash_0.x7.dcgint.t8 55.3905
R1438 flash_0.x7.dcgint.n2 flash_0.x7.dcgint.t11 55.3905
R1439 flash_0.x7.dcgint.n6 flash_0.x7.dcgint.n5 9.3005
R1440 flash_0.x7.dcgint.n5 flash_0.x7.dcgint.n4 8.9605
R1441 flash_0.x7.dcgint flash_0.x7.dcgint.n6 7.52362
R1442 flash_0.x7.dcgint.n6 flash_0.x7.dcgint.n0 1.14684
R1443 flash_0.x7.dcgint.n4 flash_0.x7.dcgint.n0 1.0086
R1444 uo_out[0].n0 uo_out[0].t0 228.901
R1445 uo_out[0].n0 uo_out[0].t1 84.4155
R1446 uo_out[0].n1 uo_out[0] 32.5825
R1447 uo_out[0].n1 uo_out[0].n0 4.88722
R1448 uo_out[0].n0 uo_out[0] 0.063
R1449 uo_out[0] uo_out[0].n1 0.016125
C0 flash_0.x4.neg_mid flash_0.x4.neg_mid_b 1.16207f
C1 flash_0.x7.VPRGPOS flash_0.x2.clkina 1.53e-19
C2 ui_in[2] flash_0.x2.stage1 5.11e-19
C3 flash_0.x7.pos_en_b flash_0.x7.vintp 0.014802f
C4 uio_in[6] uio_in[5] 0.031023f
C5 flash_0.x3.clkinb flash_0.x3.stage1 0.186066f
C6 flash_0.x7.pos_mid_b flash_0.x7.VOUT 0.781609f
C7 flash_0.x4.neg_en_b VDPWR 1.82441f
C8 flash_0.x7.VPRGNEG flash_0.x7.pos_en_b 0.22097f
C9 flash_0.x4.neg_en_b flash_0.x4.pos_mid 0.001081f
C10 flash_0.x2.clkb uo_out[0] 0.550211f
C11 flash_0.x3.stage1 flash_0.x3.clkb 0.07999f
C12 flash_0.x7.VPRGPOS flash_0.x7.pos_mid 0.417573f
C13 flash_0.x7.neg_mid flash_0.x7.VOUT 0.070044f
C14 ui_in[0] flash_0.x7.pos_mid 7.01e-20
C15 ui_in[7] ui_in[6] 0.031023f
C16 flash_0.x3.clkinb flash_0.x3.clkb 0.57785f
C17 flash_0.x7.VPRGPOS ui_in[0] 0.245007f
C18 flash_0.x4.VOUT uo_out[0] 0.031752f
C19 flash_0.x4.neg_en_b flash_0.x7.VPRGNEG 0.007732f
C20 flash_0.x2.clkb VAPWR 0.392271f
C21 flash_0.x4.pos_en_b flash_0.x7.VPRGPOS 0.064992f
C22 flash_0.x4.pos_en_b ui_in[0] 2.34221f
C23 flash_0.x7.VPRGPOS flash_0.x3.clkb 0.485638f
C24 flash_0.x7.VOUT flash_0.x7.dcgint 0.61809f
C25 flash_0.x2.clkb flash_0.x4.neg_mid_b 7.35e-19
C26 clk VAPWR 2.76692f
C27 flash_0.x7.VPRGPOS flash_0.x4.neg_mid 1.81e-19
C28 flash_0.x4.neg_mid ui_in[0] 0.003529f
C29 clk flash_0.x4.neg_mid_b 2.05e-19
C30 flash_0.x4.vintp flash_0.x4.neg_mid_b 3.34e-19
C31 flash_0.x7.VOUT ui_in[1] 0.646625f
C32 flash_0.x5.A flash_0.x7.VPRGPOS 2.9732f
C33 flash_0.x4.pos_en_b flash_0.x4.neg_mid 0.080973f
C34 flash_0.x2.clkb flash_0.x2.clkina 0.005816f
C35 flash_0.x7.neg_en_b flash_0.x7.pos_mid 0.001081f
C36 clk flash_0.x2.clkina 0.004029f
C37 flash_0.x4.neg_en_b flash_0.x4.pos_mid_b 0.013365f
C38 flash_0.x2.clka flash_0.x7.VOUT 0.01934f
C39 flash_0.x4.VOUT flash_0.x4.neg_mid_b 0.500156f
C40 flash_0.x7.neg_mid_b flash_0.x7.VOUT 0.501894f
C41 flash_0.x2.stage2 VDPWR 0.002548f
C42 flash_0.x7.neg_en_b ui_in[0] 3.05692f
C43 flash_0.x4.dcgint flash_0.x7.VOUT 0.555359f
C44 flash_0.x7.neg_mid a_20416_28577# 0.002271f
C45 clk flash_0.x3.stage1 1.05122f
C46 flash_0.x7.VOUT ui_in[2] 0.099537f
C47 a_7463_28281# VDPWR 0.08485f
C48 clk flash_0.x7.pos_mid 8.13e-22
C49 flash_0.x3.clka VAPWR 1.5347f
C50 flash_0.x2.stage2 flash_0.x7.VPRGNEG 1.79888f
C51 flash_0.x3.clkinb clk 0.350812f
C52 flash_0.x7.neg_mid uo_out[0] 0.007637f
C53 flash_0.x2.clkb flash_0.x7.VPRGPOS 0.724895f
C54 flash_0.x4.pos_mid VDPWR 0.025715f
C55 clk ui_in[0] 4.50971f
C56 flash_0.x7.VPRGPOS clk 0.234475f
C57 flash_0.x7.vintp VDPWR 0.237272f
C58 flash_0.x7.VPRGPOS flash_0.x4.vintp 0.490137f
C59 ui_in[0] flash_0.x4.vintp 8.2e-19
C60 a_20416_28577# ui_in[1] 2.08e-19
C61 a_9352_28387# a_7463_28281# 0.06129f
C62 flash_0.x7.pos_mid_b flash_0.x4.neg_mid_b 4.26e-19
C63 flash_0.x4.pos_en_b clk 3.66e-19
C64 flash_0.x2.stage2 flash_0.x3.stage2 0.035345f
C65 flash_0.x4.pos_en_b flash_0.x4.vintp 0.014802f
C66 ua[7] VDPWR 0.017072f
C67 flash_0.x4.neg_mid flash_0.x4.vintp 1.18e-20
C68 flash_0.x7.dcgint uo_out[0] 0.003294f
C69 flash_0.x5.A flash_0.x2.clkb 0.05322f
C70 a_9352_28387# VDPWR 0.04147f
C71 flash_0.x7.VPRGPOS flash_0.x4.VOUT 1.82403f
C72 ui_in[0] flash_0.x4.VOUT 0.371415f
C73 flash_0.x7.neg_mid_b a_20416_28577# 0.166835f
C74 flash_0.x5.A clk 0.00419f
C75 flash_0.x3.clka flash_0.x3.stage1 57.6093f
C76 ui_in[1] uo_out[0] 0.011391f
C77 flash_0.x7.VPRGNEG VDPWR 13.5121f
C78 flash_0.x2.stage2 flash_0.x2.clkinb 0.359889f
C79 flash_0.x4.pos_en_b flash_0.x4.VOUT 0.142413f
C80 flash_0.x4.neg_mid flash_0.x4.VOUT 0.069947f
C81 uio_in[6] uio_in[7] 0.031023f
C82 flash_0.x5.A flash_0.x4.VOUT 0.244704f
C83 flash_0.x7.neg_mid_b uo_out[0] 0.030589f
C84 flash_0.x3.clka flash_0.x3.clkinb 0.300643f
C85 a_16296_28578# uo_out[0] 0.001641f
C86 flash_0.x4.pos_mid_b VDPWR 0.302746f
C87 flash_0.x2.stage2 flash_0.x2.stage1 4.80565f
C88 flash_0.x4.pos_mid_b flash_0.x4.pos_mid 1.82667f
C89 flash_0.x4.dcgint uo_out[0] 0.002825f
C90 ui_in[1] flash_0.x4.neg_mid_b 1.66762f
C91 flash_0.x7.pos_mid_b flash_0.x7.pos_mid 1.82667f
C92 ui_in[2] uo_out[0] 2.38891f
C93 flash_0.x2.clka VAPWR 0.417222f
C94 flash_0.x7.pos_en_b flash_0.x7.VOUT 0.153015f
C95 flash_0.x3.clka flash_0.x3.clkb 1.38778f
C96 flash_0.x7.neg_mid flash_0.x7.pos_mid 4.98e-19
C97 flash_0.x7.neg_mid_b flash_0.x4.neg_mid_b 9.52e-20
C98 flash_0.x7.pos_mid_b flash_0.x7.VPRGPOS 2.35676f
C99 ua[0] VDPWR 0.053023f
C100 flash_0.x7.pos_mid_b ui_in[0] 0.126143f
C101 ui_in[7] uio_in[0] 0.031023f
C102 flash_0.x2.stage1 a_7463_28281# 1.01e-19
C103 a_16296_28578# flash_0.x4.neg_mid_b 0.166835f
C104 flash_0.x2.clka flash_0.x2.clkina 0.509107f
C105 flash_0.x4.pos_mid_b flash_0.x7.VPRGNEG 1.33e-19
C106 flash_0.x4.dcgint flash_0.x4.neg_mid_b 2.14914f
C107 flash_0.x7.neg_mid ui_in[0] 0.277486f
C108 flash_0.x7.VPRGPOS flash_0.x7.neg_mid 9.18e-20
C109 flash_0.x4.neg_en_b flash_0.x7.VOUT 0.00256f
C110 ui_in[2] flash_0.x4.neg_mid_b 0.015154f
C111 clk flash_0.x4.VOUT 0.069948f
C112 flash_0.x4.vintp flash_0.x4.VOUT 0.371874f
C113 ui_in[1] flash_0.x7.pos_mid 0.356278f
C114 flash_0.x7.VPRGPOS flash_0.x7.dcgint 4.2e-19
C115 flash_0.x7.dcgint ui_in[0] 0.146328f
C116 flash_0.x7.pos_mid_b flash_0.x7.neg_en_b 0.013365f
C117 flash_0.x7.VPRGPOS ui_in[1] 0.633798f
C118 flash_0.x7.neg_mid_b flash_0.x7.pos_mid 3.38e-20
C119 ui_in[0] ui_in[1] 8.14454f
C120 flash_0.x7.pos_en_b a_20416_28577# 3.62e-20
C121 flash_0.x7.neg_mid flash_0.x7.neg_en_b 1.5384f
C122 flash_0.x7.VPRGPOS flash_0.x2.clka 0.589813f
C123 flash_0.x4.pos_en_b ui_in[1] 0.711621f
C124 flash_0.x3.clka clk 0.013936f
C125 flash_0.x4.neg_mid ui_in[1] 0.277525f
C126 flash_0.x4.dcgint flash_0.x7.pos_mid 3.4e-19
C127 flash_0.x7.neg_mid_b ui_in[0] 1.58977f
C128 flash_0.x7.neg_mid_b flash_0.x7.VPRGPOS 0.003221f
C129 ui_in[2] flash_0.x7.pos_mid 0.017392f
C130 flash_0.x7.VPRGPOS flash_0.x6.Y 0.054645f
C131 a_16296_28578# ui_in[0] 2.08e-19
C132 flash_0.x7.pos_en_b uo_out[0] 0.01406f
C133 flash_0.x7.VPRGPOS flash_0.x4.dcgint 0.026583f
C134 flash_0.x4.dcgint ui_in[0] 0.245012f
C135 flash_0.x4.pos_en_b a_16296_28578# 3.62e-20
C136 flash_0.x5.A flash_0.x2.clka 7.82e-19
C137 flash_0.x7.neg_en_b flash_0.x7.dcgint 0.005849f
C138 flash_0.x7.pos_mid_b clk 2.14e-20
C139 flash_0.x2.stage2 flash_0.x7.VOUT 0.001251f
C140 a_16296_28578# flash_0.x4.neg_mid 0.002271f
C141 flash_0.x7.VPRGPOS ui_in[2] 0.388726f
C142 ui_in[2] ui_in[0] 0.243794f
C143 flash_0.x4.pos_en_b flash_0.x4.dcgint 0.178671f
C144 flash_0.x2.stage1 flash_0.x2.clkinb 0.189301f
C145 flash_0.x4.dcgint flash_0.x4.neg_mid 1.61e-19
C146 flash_0.x5.A flash_0.x6.Y 0.120397f
C147 flash_0.x7.neg_en_b ui_in[1] 0.031249f
C148 flash_0.x3.clkina flash_0.x3.stage2 0.20543f
C149 flash_0.x4.pos_en_b ui_in[2] 0.004173f
C150 flash_0.x7.pos_mid_b flash_0.x4.VOUT 2.87e-22
C151 flash_0.x4.neg_en_b uo_out[0] 0.00454f
C152 flash_0.x5.A ui_in[2] 0.032504f
C153 flash_0.x7.VOUT a_7463_28281# 0.128388f
C154 flash_0.x7.pos_en_b flash_0.x4.neg_mid_b 1.35e-19
C155 flash_0.x7.neg_mid_b flash_0.x7.neg_en_b 0.430883f
C156 rst_n ui_in[0] 0.031023f
C157 clk ena 0.031023f
C158 clk flash_0.x7.dcgint 2.23e-19
C159 flash_0.x7.VOUT VDPWR 2.12755f
C160 ui_in[2] flash_0.x7.neg_en_b 0.010336f
C161 flash_0.x7.VOUT flash_0.x7.vintp 0.396061f
C162 clk ui_in[1] 0.009319f
C163 uio_in[7] uo_out[0] 0.031023f
C164 flash_0.x2.clkb flash_0.x2.clka 1.38778f
C165 flash_0.x4.neg_en_b flash_0.x4.neg_mid_b 0.430883f
C166 flash_0.x2.clka clk 0.357332f
C167 flash_0.x7.VOUT a_9352_28387# 0.834577f
C168 flash_0.x7.neg_mid_b clk 9.98e-21
C169 flash_0.x4.VOUT ui_in[1] 0.456703f
C170 clk flash_0.x6.Y 0.154512f
C171 flash_0.x7.VPRGNEG flash_0.x7.VOUT 1.06096f
C172 flash_0.x2.clka flash_0.x4.VOUT 0.001465f
C173 flash_0.x7.pos_en_b flash_0.x7.pos_mid 0.595322f
C174 flash_0.x4.dcgint flash_0.x4.vintp 1.54e-20
C175 clk ui_in[2] 2.12761f
C176 flash_0.x2.stage2 uo_out[0] 0.002424f
C177 flash_0.x6.Y flash_0.x4.VOUT 0.044456f
C178 ui_in[2] flash_0.x4.vintp 0.00728f
C179 flash_0.x7.pos_mid_b flash_0.x7.neg_mid 0.001246f
C180 a_16296_28578# flash_0.x4.VOUT 0.017698f
C181 flash_0.x7.VPRGPOS flash_0.x7.pos_en_b 0.077604f
C182 flash_0.x7.pos_en_b ui_in[0] 0.712549f
C183 flash_0.x4.pos_mid_b flash_0.x7.VOUT 5.14e-19
C184 flash_0.x4.dcgint flash_0.x4.VOUT 0.619301f
C185 ui_in[2] flash_0.x4.VOUT 0.226315f
C186 a_20416_28577# VDPWR 0.106135f
C187 rst_n clk 0.031023f
C188 ui_in[3] ui_in[2] 0.031023f
C189 flash_0.x7.pos_mid_b flash_0.x7.dcgint 0.009409f
C190 flash_0.x2.stage2 VAPWR 7.897181f
C191 ui_in[4] ui_in[5] 0.031023f
C192 flash_0.x2.stage2 flash_0.x4.neg_mid_b 0.002851f
C193 flash_0.x4.neg_en_b flash_0.x7.VPRGPOS 0.002081f
C194 flash_0.x4.neg_en_b ui_in[0] 0.030971f
C195 flash_0.x7.pos_mid_b ui_in[1] 0.774227f
C196 uo_out[0] VDPWR 0.609895f
C197 flash_0.x7.neg_mid flash_0.x7.dcgint 1.61e-19
C198 flash_0.x4.pos_en_b flash_0.x4.neg_en_b 0.337454f
C199 flash_0.x2.stage2 flash_0.x2.clkina 0.206461f
C200 uio_in[1] uio_in[0] 0.031023f
C201 flash_0.x7.pos_en_b flash_0.x7.neg_en_b 0.337454f
C202 flash_0.x4.neg_en_b flash_0.x4.neg_mid 1.5384f
C203 flash_0.x7.VOUT flash_0.x2.stage1 0.001452f
C204 flash_0.x7.VPRGNEG a_20416_28577# 0.062489f
C205 flash_0.x7.neg_mid ui_in[1] 0.003547f
C206 flash_0.x7.neg_mid_b flash_0.x7.pos_mid_b 0.428431f
C207 uio_in[5] uio_in[4] 0.031023f
C208 flash_0.x7.pos_mid_b flash_0.x4.dcgint 4.14e-19
C209 flash_0.x7.neg_mid_b flash_0.x7.neg_mid 1.16207f
C210 VAPWR VDPWR 0.724319f
C211 flash_0.x7.VPRGNEG uo_out[0] 3.06829f
C212 VDPWR flash_0.x4.neg_mid_b 1.912801f
C213 flash_0.x7.pos_mid_b ui_in[2] 0.039178f
C214 flash_0.x4.pos_mid flash_0.x4.neg_mid_b 3.38e-20
C215 flash_0.x7.dcgint ui_in[1] 0.239891f
C216 flash_0.x7.pos_en_b clk 1.99e-20
C217 flash_0.x7.neg_mid ui_in[2] 0.001615f
C218 flash_0.x7.neg_mid_b flash_0.x7.dcgint 2.14914f
C219 flash_0.x3.stage2 uo_out[0] 0.080392f
C220 flash_0.x2.stage2 flash_0.x7.VPRGPOS 0.757314f
C221 flash_0.x7.VPRGNEG VAPWR 2.20506f
C222 flash_0.x7.neg_mid_b ui_in[1] 0.208234f
C223 flash_0.x7.VPRGNEG flash_0.x4.neg_mid_b 2.19355f
C224 flash_0.x2.stage2 flash_0.x3.clkb 4.24817f
C225 ui_in[2] flash_0.x7.dcgint 0.039612f
C226 flash_0.x4.dcgint ui_in[1] 0.278517f
C227 flash_0.x5.A flash_0.x2.stage2 0.002905f
C228 flash_0.x7.pos_mid VDPWR 0.018345f
C229 ui_in[2] ui_in[1] 4.33478f
C230 VAPWR flash_0.x3.stage2 1.42027f
C231 flash_0.x7.VPRGPOS a_7463_28281# 0.169831f
C232 flash_0.x4.pos_mid_b flash_0.x4.neg_mid_b 0.428431f
C233 flash_0.x7.vintp flash_0.x7.pos_mid 0.007513f
C234 flash_0.x2.clka ui_in[2] 0.003846f
C235 flash_0.x7.neg_mid_b flash_0.x4.dcgint 1.52e-19
C236 flash_0.x4.neg_en_b flash_0.x4.VOUT 0.293379f
C237 flash_0.x7.VPRGPOS VDPWR 3.63662f
C238 ui_in[0] VDPWR 3.543282f
C239 flash_0.x7.neg_mid_b ui_in[2] 0.034018f
C240 flash_0.x7.VPRGPOS flash_0.x4.pos_mid 0.416622f
C241 VAPWR flash_0.x2.clkinb 1.65827f
C242 ui_in[0] flash_0.x4.pos_mid 0.343817f
C243 ui_in[2] flash_0.x6.Y 0.447688f
C244 flash_0.x7.VPRGPOS flash_0.x7.vintp 0.490248f
C245 flash_0.x4.pos_en_b VDPWR 1.861514f
C246 flash_0.x4.pos_en_b flash_0.x4.pos_mid 0.595322f
C247 flash_0.x4.neg_mid VDPWR 1.39258f
C248 flash_0.x4.dcgint ui_in[2] 0.014403f
C249 ui_in[3] ui_in[4] 0.031023f
C250 flash_0.x4.neg_mid flash_0.x4.pos_mid 4.98e-19
C251 uio_in[3] uio_in[2] 0.031023f
C252 flash_0.x2.clkina flash_0.x2.clkinb 0.886684f
C253 flash_0.x5.A VDPWR 2.1939f
C254 flash_0.x7.pos_mid_b flash_0.x7.pos_en_b 0.391527f
C255 flash_0.x3.stage1 flash_0.x3.stage2 5.8896f
C256 flash_0.x7.VPRGPOS a_9352_28387# 0.393793f
C257 VAPWR flash_0.x2.stage1 5.931509f
C258 flash_0.x7.VPRGPOS flash_0.x7.VPRGNEG 1.33754f
C259 flash_0.x7.VPRGNEG ui_in[0] 0.063928f
C260 flash_0.x7.neg_mid flash_0.x7.pos_en_b 0.080973f
C261 flash_0.x2.stage2 flash_0.x2.clkb 58.9902f
C262 uio_in[2] uio_in[1] 0.031023f
C263 flash_0.x7.neg_en_b VDPWR 1.678f
C264 flash_0.x4.pos_en_b flash_0.x7.VPRGNEG 0.232602f
C265 flash_0.x2.clkina flash_0.x2.stage1 0.01805f
C266 flash_0.x3.clkinb flash_0.x3.stage2 0.358189f
C267 flash_0.x4.neg_mid flash_0.x7.VPRGNEG 0.976831f
C268 flash_0.x5.A a_9352_28387# 0.868312f
C269 flash_0.x3.clkina VAPWR 1.05609f
C270 flash_0.x4.pos_mid_b ui_in[0] 0.762651f
C271 flash_0.x7.VPRGPOS flash_0.x3.stage2 1.93468f
C272 flash_0.x4.pos_mid_b flash_0.x7.VPRGPOS 2.26733f
C273 flash_0.x7.pos_en_b flash_0.x7.dcgint 0.178671f
C274 flash_0.x4.pos_en_b flash_0.x4.pos_mid_b 0.391527f
C275 flash_0.x3.clkb flash_0.x3.stage2 59.0307f
C276 flash_0.x3.stage1 flash_0.x2.stage1 0.030249f
C277 flash_0.x4.pos_mid_b flash_0.x4.neg_mid 0.001246f
C278 flash_0.x7.VPRGNEG flash_0.x7.neg_en_b 0.007055f
C279 flash_0.x7.VPRGPOS flash_0.x2.clkinb 2.41e-19
C280 flash_0.x7.pos_en_b ui_in[1] 2.34386f
C281 flash_0.x2.clkb VDPWR 0.024098f
C282 flash_0.x7.VPRGPOS ua[0] 0.043554f
C283 flash_0.x7.VOUT a_20416_28577# 0.017698f
C284 clk VDPWR 0.461416f
C285 flash_0.x4.vintp VDPWR 0.237277f
C286 clk flash_0.x4.pos_mid 1.68e-20
C287 flash_0.x4.VOUT a_7463_28281# 0.069775f
C288 flash_0.x4.vintp flash_0.x4.pos_mid 0.007513f
C289 flash_0.x3.clkina flash_0.x3.stage1 0.013783f
C290 flash_0.x7.neg_mid_b flash_0.x7.pos_en_b 0.743046f
C291 flash_0.x7.VPRGPOS flash_0.x2.stage1 0.125764f
C292 flash_0.x2.stage2 flash_0.x3.clka 0.011129f
C293 flash_0.x4.VOUT VDPWR 2.542964f
C294 flash_0.x4.neg_en_b ui_in[1] 3.07359f
C295 flash_0.x4.dcgint flash_0.x7.pos_en_b 1.62e-19
C296 flash_0.x2.clkb a_9352_28387# 0.002716f
C297 flash_0.x7.VOUT uo_out[0] 0.093374f
C298 flash_0.x4.VOUT flash_0.x4.pos_mid 0.013006f
C299 flash_0.x3.clkb flash_0.x2.stage1 7.28e-19
C300 flash_0.x3.clkina flash_0.x3.clkinb 0.886684f
C301 flash_0.x2.clkb flash_0.x7.VPRGNEG 0.572269f
C302 flash_0.x7.pos_en_b ui_in[2] 0.007039f
C303 ui_in[5] ui_in[6] 0.031023f
C304 flash_0.x4.neg_en_b a_16296_28578# 6.87e-21
C305 a_9352_28387# flash_0.x4.VOUT 0.039663f
C306 flash_0.x3.clkina flash_0.x3.clkb 0.005939f
C307 flash_0.x4.neg_en_b flash_0.x4.dcgint 0.005849f
C308 flash_0.x7.VPRGNEG flash_0.x4.VOUT 0.387788f
C309 uio_in[3] uio_in[4] 0.031023f
C310 flash_0.x7.VOUT flash_0.x4.neg_mid_b 0.002509f
C311 flash_0.x4.pos_mid_b clk 5.23e-19
C312 flash_0.x4.neg_en_b ui_in[2] 0.001238f
C313 flash_0.x4.pos_mid_b flash_0.x4.vintp 0.252393f
C314 flash_0.x2.clkb flash_0.x2.clkinb 0.577668f
C315 clk flash_0.x2.clkinb 0.350812f
C316 flash_0.x4.pos_mid_b flash_0.x4.VOUT 0.256021f
C317 flash_0.x7.pos_mid_b VDPWR 0.286404f
C318 ua[0] clk 0.304224f
C319 flash_0.x7.pos_mid_b flash_0.x7.vintp 0.252393f
C320 a_20416_28577# uo_out[0] 0.001639f
C321 flash_0.x7.neg_mid VDPWR 1.38354f
C322 flash_0.x2.clkb flash_0.x2.stage1 0.080777f
C323 flash_0.x2.stage2 flash_0.x2.clka 1.79536f
C324 clk flash_0.x2.stage1 2.76362f
C325 flash_0.x7.neg_mid flash_0.x7.vintp 1.18e-20
C326 flash_0.x7.VOUT flash_0.x7.pos_mid 0.349932f
C327 flash_0.x7.pos_mid_b flash_0.x7.VPRGNEG 1.33e-19
C328 flash_0.x3.clka flash_0.x3.stage2 1.79536f
C329 flash_0.x7.dcgint VDPWR 0.007589f
C330 flash_0.x4.VOUT flash_0.x2.stage1 3.9e-20
C331 flash_0.x3.clkina clk 0.004029f
C332 flash_0.x2.clka a_7463_28281# 0.011214f
C333 flash_0.x7.neg_mid flash_0.x7.VPRGNEG 0.976831f
C334 flash_0.x7.VPRGPOS flash_0.x7.VOUT 4.05971f
C335 flash_0.x7.VOUT ui_in[0] 0.473707f
C336 flash_0.x7.vintp flash_0.x7.dcgint 1.54e-20
C337 ui_in[1] VDPWR 3.657281f
C338 flash_0.x4.pos_en_b flash_0.x7.VOUT 0.023223f
C339 flash_0.x7.vintp ui_in[1] 0.006255f
C340 flash_0.x4.neg_mid flash_0.x7.VOUT 1.16e-19
C341 flash_0.x7.neg_mid_b VDPWR 1.799591f
C342 uo_out[0] flash_0.x4.neg_mid_b 0.030267f
C343 flash_0.x5.A flash_0.x7.VOUT 0.207778f
C344 flash_0.x6.Y VDPWR 7.946081f
C345 a_16296_28578# VDPWR 0.106132f
C346 flash_0.x4.neg_en_b flash_0.x7.pos_en_b 0.005326f
C347 ui_in[2] a_7463_28281# 0.196624f
C348 flash_0.x7.neg_mid_b flash_0.x7.vintp 3.34e-19
C349 flash_0.x3.clka flash_0.x2.stage1 4.27357f
C350 flash_0.x4.dcgint VDPWR 0.047507f
C351 flash_0.x7.VPRGNEG ui_in[1] 0.065673f
C352 flash_0.x2.clka a_9352_28387# 0.002596f
C353 ui_in[2] VDPWR 3.521599f
C354 flash_0.x7.VOUT flash_0.x7.neg_en_b 0.293369f
C355 ui_in[2] flash_0.x4.pos_mid 0.022101f
C356 ui_in[2] flash_0.x7.vintp 0.007287f
C357 flash_0.x7.neg_mid_b flash_0.x7.VPRGNEG 2.18563f
C358 flash_0.x3.clka flash_0.x3.clkina 0.509107f
C359 a_16296_28578# flash_0.x7.VPRGNEG 0.062517f
C360 flash_0.x4.pos_mid_b ui_in[1] 0.022428f
C361 flash_0.x2.clkina VAPWR 1.04794f
C362 flash_0.x4.dcgint flash_0.x7.VPRGNEG 4.72e-19
C363 flash_0.x2.clkb flash_0.x7.VOUT 0.084343f
C364 flash_0.x7.VOUT clk 2.11e-20
C365 flash_0.x2.clka flash_0.x2.clkinb 0.30061f
C366 flash_0.x3.stage1 VAPWR 4.90996f
C367 ui_in[0] uo_out[0] 0.016476f
C368 flash_0.x4.pos_mid_b flash_0.x4.dcgint 0.009409f
C369 flash_0.x7.VPRGPOS uo_out[0] 2.61882f
C370 flash_0.x4.pos_mid_b ui_in[2] 0.047751f
C371 flash_0.x4.pos_en_b uo_out[0] 0.012717f
C372 flash_0.x4.neg_mid uo_out[0] 0.007647f
C373 flash_0.x7.VOUT flash_0.x4.VOUT 0.38054f
C374 flash_0.x7.pos_mid flash_0.x4.neg_mid_b 0.001667f
C375 ua[0] flash_0.x6.Y 0.290173f
C376 flash_0.x3.clkinb VAPWR 1.66476f
C377 flash_0.x2.clka flash_0.x2.stage1 57.610302f
C378 flash_0.x7.neg_en_b a_20416_28577# 6.87e-21
C379 flash_0.x5.A uo_out[0] 0.225691f
C380 ui_in[0] flash_0.x4.neg_mid_b 0.209459f
C381 flash_0.x7.VPRGPOS flash_0.x4.neg_mid_b 0.008594f
C382 ua[0] ui_in[2] 0.009579f
C383 VAPWR flash_0.x3.clkb 0.370933f
C384 flash_0.x4.pos_en_b flash_0.x4.neg_mid_b 0.743046f
C385 flash_0.x7.neg_en_b uo_out[0] 0.00488f
C386 flash_0.x7.pos_en_b VDPWR 1.804284f
C387 ua[1] VGND 0.146962f
C388 ua[2] VGND 0.146962f
C389 ua[3] VGND 0.146962f
C390 ua[4] VGND 0.146962f
C391 ua[5] VGND 0.146962f
C392 ua[6] VGND 0.146962f
C393 ua[7] VGND 0.128006f
C394 ena VGND 0.070385f
C395 rst_n VGND 0.042875f
C396 ui_in[3] VGND 0.042875f
C397 ui_in[4] VGND 0.042875f
C398 ui_in[5] VGND 0.042875f
C399 ui_in[6] VGND 0.042875f
C400 ui_in[7] VGND 0.042875f
C401 uio_in[0] VGND 0.042875f
C402 uio_in[1] VGND 0.042875f
C403 uio_in[2] VGND 0.042875f
C404 uio_in[3] VGND 0.042875f
C405 uio_in[4] VGND 0.042875f
C406 uio_in[5] VGND 0.042875f
C407 uio_in[6] VGND 0.042875f
C408 uio_in[7] VGND 0.042875f
C409 ui_in[0] VGND 23.129925f
C410 ui_in[1] VGND 20.58311f
C411 uo_out[0] VGND 13.615086f
C412 ui_in[2] VGND 15.773119f
C413 clk VGND 25.498606f
C414 ua[0] VGND 35.369205f
C415 VDPWR VGND 98.75901f
C416 VAPWR VGND 43.180836f
C417 flash_0.x7.vintp VGND 0.039625f
C418 flash_0.x4.vintp VGND 0.051188f
C419 flash_0.x7.pos_mid VGND 1.29059f
C420 flash_0.x7.pos_mid_b VGND 3.938035f
C421 flash_0.x4.pos_mid VGND 1.31994f
C422 flash_0.x4.pos_mid_b VGND 3.985879f
C423 flash_0.x6.Y VGND 13.6985f
C424 flash_0.x7.neg_en_b VGND 3.319393f
C425 flash_0.x7.neg_mid VGND 0.210934f
C426 a_20416_28577# VGND 0.048706f
C427 flash_0.x7.neg_mid_b VGND 4.319581f
C428 flash_0.x7.pos_en_b VGND 7.747194f
C429 flash_0.x4.neg_en_b VGND 3.199902f
C430 flash_0.x4.neg_mid VGND 0.206959f
C431 a_16296_28578# VGND 0.047639f
C432 flash_0.x4.neg_mid_b VGND 4.854208f
C433 flash_0.x4.pos_en_b VGND 7.770404f
C434 a_9352_28387# VGND 0.21567f
C435 flash_0.x4.VOUT VGND 6.814736f
C436 a_7463_28281# VGND 0.801294f
C437 flash_0.x2.clkb VGND 63.13064f
C438 flash_0.x2.clka VGND 62.52466f
C439 flash_0.x2.clkinb VGND 3.11026f
C440 flash_0.x2.clkina VGND 1.57797f
C441 flash_0.x3.clkb VGND 66.16767f
C442 flash_0.x3.clka VGND 65.171394f
C443 flash_0.x3.clkinb VGND 3.10612f
C444 flash_0.x3.clkina VGND 1.5755f
C445 flash_0.x7.dcgint VGND 3.309877f
C446 flash_0.x4.dcgint VGND 2.988657f
C447 flash_0.x5.A VGND 5.742692f
C448 flash_0.x7.VOUT VGND 12.457275f
C449 flash_0.x7.VPRGNEG VGND 80.182205f
C450 flash_0.x2.stage2 VGND 15.4695f
C451 flash_0.x2.stage1 VGND 18.413f
C452 flash_0.x7.VPRGPOS VGND 0.148564p
C453 flash_0.x3.stage2 VGND 24.3058f
C454 flash_0.x3.stage1 VGND 23.173801f
C455 uo_out[0].t0 VGND 0.038292f
C456 uo_out[0].t1 VGND 0.037022f
C457 uo_out[0].n0 VGND 0.257992f
C458 uo_out[0].n1 VGND 3.39873f
C459 flash_0.x7.dcgint.t0 VGND 0.016015f
C460 flash_0.x7.dcgint.t1 VGND 0.016015f
C461 flash_0.x7.dcgint.t2 VGND 0.016015f
C462 flash_0.x7.dcgint.t7 VGND 0.017561f
C463 flash_0.x7.dcgint.n0 VGND 0.05401f
C464 flash_0.x7.dcgint.t4 VGND 0.017266f
C465 flash_0.x7.dcgint.t9 VGND 0.355987f
C466 flash_0.x7.dcgint.t5 VGND 0.222316f
C467 flash_0.x7.dcgint.t3 VGND 0.280884f
C468 flash_0.x7.dcgint.t6 VGND 0.004616f
C469 flash_0.x7.dcgint.t10 VGND 0.004616f
C470 flash_0.x7.dcgint.n1 VGND 0.009325f
C471 flash_0.x7.dcgint.t8 VGND 0.004616f
C472 flash_0.x7.dcgint.t11 VGND 0.004616f
C473 flash_0.x7.dcgint.n2 VGND 0.009325f
C474 flash_0.x7.dcgint.n3 VGND 0.045712f
C475 flash_0.x7.dcgint.n4 VGND 0.233815f
C476 flash_0.x7.dcgint.n5 VGND 0.046322f
C477 flash_0.x7.dcgint.n6 VGND 0.34091f
C478 flash_0.x2.clka.t0 VGND 0.011299f
C479 flash_0.x2.clka.t1 VGND 0.017732f
C480 ui_in[2].t2 VGND 0.727097f
C481 ui_in[2].t0 VGND 0.69579f
C482 ui_in[2].n0 VGND 0.550323f
C483 ui_in[2].t1 VGND 0.186184f
C484 ui_in[2].n1 VGND 1.11593f
C485 ui_in[2].n2 VGND 4.46526f
C486 flash_0.x4.pos_en_b.n0 VGND 0.032452f
C487 flash_0.x4.pos_en_b.n1 VGND 0.766491f
C488 flash_0.x4.pos_en_b.t4 VGND 0.932199f
C489 flash_0.x4.pos_en_b.t5 VGND 0.216253f
C490 flash_0.x4.pos_en_b.t6 VGND 0.216253f
C491 flash_0.x4.pos_en_b.t1 VGND 0.010089f
C492 flash_0.x4.pos_en_b.t0 VGND 0.010089f
C493 flash_0.x4.pos_en_b.t2 VGND 0.008975f
C494 flash_0.x4.pos_en_b.t3 VGND 0.008975f
C495 flash_0.x3.clkb.t0 VGND 0.012451f
C496 flash_0.x3.clkb.t1 VGND 0.01954f
C497 flash_0.x3.clka.t0 VGND 0.012142f
C498 flash_0.x3.clka.t1 VGND 0.019055f
C499 w_7728_24730.t2 VGND 6.5007f
C500 w_7728_24730.t0 VGND 6.37557f
C501 w_7728_24730.t1 VGND 0.011863f
C502 w_7728_24730.t3 VGND 0.01187f
C503 flash_0.x7.VOUT.n0 VGND 2.03422f
C504 flash_0.x7.VOUT.n1 VGND 0.036039f
C505 flash_0.x7.VOUT.t11 VGND 0.015115f
C506 flash_0.x7.VOUT.t13 VGND 0.003984f
C507 flash_0.x7.VOUT.t10 VGND 0.003984f
C508 flash_0.x7.VOUT.n2 VGND 0.008188f
C509 flash_0.x7.VOUT.t8 VGND 0.003984f
C510 flash_0.x7.VOUT.t9 VGND 0.003984f
C511 flash_0.x7.VOUT.n3 VGND 0.008184f
C512 flash_0.x7.VOUT.t12 VGND 0.015115f
C513 flash_0.x7.VOUT.t0 VGND 0.013679f
C514 flash_0.x7.VOUT.t1 VGND 0.013673f
C515 flash_0.x7.VOUT.n4 VGND 0.034644f
C516 flash_0.x7.VOUT.n5 VGND 0.035068f
C517 flash_0.x7.VOUT.n6 VGND 0.034644f
C518 flash_0.x7.VOUT.n7 VGND 0.025905f
C519 flash_0.x7.VOUT.n8 VGND 0.224312f
C520 flash_0.x7.VOUT.t14 VGND 0.282327f
C521 flash_0.x7.VOUT.n11 VGND 0.224312f
C522 flash_0.x7.VOUT.n12 VGND 0.025537f
C523 flash_0.x7.VOUT.t7 VGND 0.01411f
C524 flash_0.x7.VOUT.t5 VGND 0.01411f
C525 flash_0.x7.VOUT.t6 VGND 0.003984f
C526 flash_0.x7.VOUT.t4 VGND 0.003984f
C527 flash_0.x7.VOUT.n13 VGND 0.008184f
C528 flash_0.x7.VOUT.t2 VGND 0.003984f
C529 flash_0.x7.VOUT.t3 VGND 0.003984f
C530 flash_0.x7.VOUT.n14 VGND 0.008184f
C531 ui_in[0].t6 VGND 0.037781f
C532 ui_in[0].n0 VGND 0.057717f
C533 ui_in[0].t14 VGND 0.037781f
C534 ui_in[0].n1 VGND 0.14905f
C535 ui_in[0].t8 VGND 0.037781f
C536 ui_in[0].n2 VGND 0.109725f
C537 ui_in[0].t9 VGND 0.037781f
C538 ui_in[0].n3 VGND 0.14905f
C539 ui_in[0].t0 VGND 0.037781f
C540 ui_in[0].n4 VGND 0.057717f
C541 ui_in[0].t10 VGND 0.037781f
C542 ui_in[0].n5 VGND 0.146838f
C543 ui_in[0].n6 VGND 0.408027f
C544 ui_in[0].t16 VGND 0.266104f
C545 ui_in[0].t12 VGND 0.278064f
C546 ui_in[0].n7 VGND 0.44849f
C547 ui_in[0].n8 VGND 0.330488f
C548 ui_in[0].t5 VGND 0.266104f
C549 ui_in[0].t2 VGND 0.278064f
C550 ui_in[0].n9 VGND 0.44849f
C551 ui_in[0].n10 VGND 0.227519f
C552 ui_in[0].n11 VGND 0.226122f
C553 ui_in[0].n12 VGND 0.127227f
C554 ui_in[0].n13 VGND 1.01912f
C555 ui_in[0].t3 VGND 0.22275f
C556 ui_in[0].t1 VGND 0.20481f
C557 ui_in[0].n14 VGND 0.313943f
C558 ui_in[0].n15 VGND 0.120049f
C559 ui_in[0].n16 VGND 0.1624f
C560 ui_in[0].t7 VGND 0.266104f
C561 ui_in[0].t4 VGND 0.278064f
C562 ui_in[0].n17 VGND 0.44849f
C563 ui_in[0].n18 VGND 0.223258f
C564 ui_in[0].n19 VGND 0.099266f
C565 ui_in[0].t17 VGND 0.266104f
C566 ui_in[0].t15 VGND 0.278064f
C567 ui_in[0].n20 VGND 0.44849f
C568 ui_in[0].n21 VGND 0.223258f
C569 ui_in[0].n22 VGND 0.099844f
C570 ui_in[0].n23 VGND 0.313671f
C571 ui_in[0].t13 VGND 0.22275f
C572 ui_in[0].t11 VGND 0.20481f
C573 ui_in[0].n24 VGND 0.313943f
C574 ui_in[0].n25 VGND 0.129255f
C575 ui_in[0].n26 VGND 0.508238f
C576 ui_in[0].n27 VGND 3.80721f
C577 flash_0.x5.A.n0 VGND 0.493086f
C578 flash_0.x5.A.n1 VGND 0.103919f
C579 flash_0.x5.A.t5 VGND 0.417187f
C580 flash_0.x5.A.t4 VGND 0.436255f
C581 flash_0.x5.A.t0 VGND 0.014943f
C582 flash_0.x5.A.n2 VGND 0.065317f
C583 flash_0.x5.A.n3 VGND 0.639596f
C584 flash_0.x5.A.n4 VGND 0.639596f
C585 flash_0.x5.A.n5 VGND 0.068344f
C586 flash_0.x5.A.n6 VGND 0.114375f
C587 flash_0.x5.A.t2 VGND 0.747064f
C588 flash_0.x5.A.n9 VGND 0.114375f
C589 flash_0.x5.A.n10 VGND 0.06833f
C590 flash_0.x5.A.t3 VGND 0.110389f
C591 flash_0.x5.A.t1 VGND 0.169707f
C592 flash_0.x5.A.n11 VGND 0.595547f
C593 flash_0.x6.Y.t0 VGND 0.038013f
C594 flash_0.x7.neg_mid_b.n0 VGND 0.539196f
C595 flash_0.x7.neg_mid_b.t10 VGND 0.243062f
C596 flash_0.x7.neg_mid_b.t9 VGND 0.243062f
C597 flash_0.x7.neg_mid_b.n1 VGND 0.341911f
C598 flash_0.x7.neg_mid_b.n2 VGND 0.140489f
C599 flash_0.x7.neg_mid_b.t0 VGND 0.027096f
C600 flash_0.x7.neg_mid_b.t3 VGND 0.007678f
C601 flash_0.x7.neg_mid_b.t1 VGND 0.007678f
C602 flash_0.x7.neg_mid_b.n3 VGND 0.015666f
C603 flash_0.x7.neg_mid_b.t15 VGND 0.085863f
C604 flash_0.x7.neg_mid_b.t6 VGND 0.02816f
C605 flash_0.x7.neg_mid_b.t7 VGND 0.067252f
C606 flash_0.x7.neg_mid_b.t8 VGND 0.122491f
C607 flash_0.x7.neg_mid_b.t11 VGND 0.067252f
C608 flash_0.x7.neg_mid_b.t13 VGND 0.122491f
C609 flash_0.x7.neg_mid_b.t12 VGND 0.067252f
C610 flash_0.x7.neg_mid_b.t14 VGND 0.122491f
C611 flash_0.x7.neg_mid_b.t4 VGND 0.007678f
C612 flash_0.x7.neg_mid_b.t2 VGND 0.007678f
C613 flash_0.x7.neg_mid_b.n4 VGND 0.015661f
C614 flash_0.x7.neg_mid_b.t5 VGND 0.02709f
C615 flash_0.x7.neg_en_b.t2 VGND 0.038945f
C616 flash_0.x7.neg_en_b.t9 VGND 0.052338f
C617 flash_0.x7.neg_en_b.t5 VGND 0.051225f
C618 flash_0.x7.neg_en_b.t7 VGND 0.051225f
C619 flash_0.x7.neg_en_b.t4 VGND 0.051225f
C620 flash_0.x7.neg_en_b.t8 VGND 0.051201f
C621 flash_0.x7.neg_en_b.t6 VGND 0.051201f
C622 flash_0.x7.neg_en_b.t1 VGND 0.036466f
C623 flash_0.x7.neg_en_b.t3 VGND 0.032439f
C624 flash_0.x7.neg_en_b.t0 VGND 0.032439f
C625 ua[0].t3 VGND 0.00285f
C626 ua[0].t2 VGND 0.716764f
C627 ua[0].n0 VGND 0.259475f
C628 ua[0].t1 VGND 0.002851f
C629 ua[0].n1 VGND 0.024193f
C630 ua[0].n2 VGND 0.02427f
C631 ua[0].n4 VGND 0.042071f
C632 ua[0].n5 VGND 0.02521f
C633 ua[0].n6 VGND 0.281781f
C634 ua[0].t0 VGND 0.430674f
C635 ua[0].n8 VGND 0.042071f
C636 ua[0].n9 VGND 0.281781f
C637 ua[0].n10 VGND 0.015559f
C638 ua[0].n11 VGND 0.0156f
C639 ua[0].n12 VGND -0.00395f
C640 ua[0].n13 VGND 0.015585f
C641 ua[0].n14 VGND 1.92631f
C642 VDPWR.t41 VGND 0.004533f
C643 VDPWR.t38 VGND 0.004533f
C644 VDPWR.n0 VGND 0.009293f
C645 VDPWR.t7 VGND 0.001565f
C646 VDPWR.t56 VGND 0.001565f
C647 VDPWR.n1 VGND 0.00313f
C648 VDPWR.n2 VGND 0.004476f
C649 VDPWR.t11 VGND 0.001565f
C650 VDPWR.t28 VGND 0.001565f
C651 VDPWR.n3 VGND 0.00313f
C652 VDPWR.n4 VGND 0.004476f
C653 VDPWR.n5 VGND 0.094814f
C654 VDPWR.t3 VGND 0.001565f
C655 VDPWR.t52 VGND 0.001565f
C656 VDPWR.n6 VGND 0.00313f
C657 VDPWR.n7 VGND 0.004476f
C658 VDPWR.t8 VGND 0.001565f
C659 VDPWR.t55 VGND 0.001565f
C660 VDPWR.n8 VGND 0.00313f
C661 VDPWR.n9 VGND 0.004476f
C662 VDPWR.n10 VGND 0.146582f
C663 VDPWR.t24 VGND 0.001565f
C664 VDPWR.t57 VGND 0.001565f
C665 VDPWR.n11 VGND 0.00313f
C666 VDPWR.n12 VGND 0.004476f
C667 VDPWR.t10 VGND 0.001565f
C668 VDPWR.t48 VGND 0.001565f
C669 VDPWR.n13 VGND 0.00313f
C670 VDPWR.n14 VGND 0.004476f
C671 VDPWR.n15 VGND 0.030697f
C672 VDPWR.n16 VGND 0.092993f
C673 VDPWR.t50 VGND 0.004533f
C674 VDPWR.t26 VGND 0.004533f
C675 VDPWR.n17 VGND 0.009293f
C676 VDPWR.n18 VGND 0.025631f
C677 VDPWR.n19 VGND 0.058575f
C678 VDPWR.n20 VGND 12.4768f
C679 VDPWR.n21 VGND 0.047001f
C680 VDPWR.t46 VGND 0.00592f
C681 VDPWR.n22 VGND 0.087115f
C682 VDPWR.n23 VGND 0.087207f
C683 VDPWR.n25 VGND 0.149716f
C684 VDPWR.n26 VGND 0.089131f
C685 VDPWR.n27 VGND 1.02311f
C686 VDPWR.t45 VGND 1.64207f
C687 VDPWR.n29 VGND 0.149716f
C688 VDPWR.n30 VGND 1.02311f
C689 VDPWR.n31 VGND 0.048652f
C690 VDPWR.n32 VGND 0.048666f
C691 VDPWR.n33 VGND 0.370974f
C692 VDPWR.t54 VGND 0.011501f
C693 VDPWR.n34 VGND 0.027153f
C694 VDPWR.n35 VGND 0.002716f
C695 VDPWR.n36 VGND 0.026195f
C696 VDPWR.n37 VGND 0.20679f
C697 VDPWR.n38 VGND 0.20679f
C698 VDPWR.n39 VGND 0.013213f
C699 VDPWR.n40 VGND 0.02444f
C700 VDPWR.n41 VGND 0.025845f
C701 VDPWR.t53 VGND 0.321959f
C702 VDPWR.n44 VGND 0.025845f
C703 VDPWR.n45 VGND 0.02444f
C704 VDPWR.n46 VGND 0.013174f
C705 VDPWR.n47 VGND 0.038779f
C706 VDPWR.n48 VGND 0.45602f
C707 VDPWR.n49 VGND 0.14638f
C708 VDPWR.n50 VGND 1.04504f
C709 VDPWR.t5 VGND 0.011501f
C710 VDPWR.n51 VGND 0.027153f
C711 VDPWR.n52 VGND 0.002716f
C712 VDPWR.n53 VGND 0.026195f
C713 VDPWR.n54 VGND 0.20679f
C714 VDPWR.n55 VGND 0.20679f
C715 VDPWR.n56 VGND 0.013213f
C716 VDPWR.n57 VGND 0.02444f
C717 VDPWR.n58 VGND 0.025845f
C718 VDPWR.t4 VGND 0.321959f
C719 VDPWR.n61 VGND 0.025845f
C720 VDPWR.n62 VGND 0.02444f
C721 VDPWR.n63 VGND 0.013174f
C722 VDPWR.n64 VGND 0.095248f
C723 VDPWR.n65 VGND 1.55096f
C724 VDPWR.t1 VGND 0.004533f
C725 VDPWR.t30 VGND 0.004533f
C726 VDPWR.n66 VGND 0.009293f
C727 VDPWR.n67 VGND 0.076846f
C728 VDPWR.n68 VGND 0.024591f
C729 VDPWR.n69 VGND 0.054924f
C730 VDPWR.n70 VGND 0.061618f
C731 VDPWR.n71 VGND 0.061618f
C732 VDPWR.n72 VGND 0.478933f
C733 VDPWR.t22 VGND 0.190001f
C734 VDPWR.t14 VGND 0.132715f
C735 VDPWR.t32 VGND 0.074358f
C736 VDPWR.t16 VGND 0.090359f
C737 VDPWR.t12 VGND 0.148716f
C738 VDPWR.t18 VGND 0.148716f
C739 VDPWR.t20 VGND 0.192013f
C740 VDPWR.t59 VGND 0.049545f
C741 VDPWR.t58 VGND 0.049545f
C742 VDPWR.n73 VGND 0.068002f
C743 VDPWR.n74 VGND 0.01319f
C744 VDPWR.n75 VGND 0.049068f
C745 VDPWR.n76 VGND 0.057729f
C746 VDPWR.n77 VGND 0.055525f
C747 VDPWR.n78 VGND 0.027565f
C748 VDPWR.n79 VGND 0.061913f
C749 VDPWR.n80 VGND 0.259805f
C750 VDPWR.n81 VGND 0.125237f
C751 VDPWR.t42 VGND 0.270154f
C752 VDPWR.t0 VGND 0.21587f
C753 VDPWR.n82 VGND 0.186521f
C754 VDPWR.t29 VGND 0.37276f
C755 VDPWR.n83 VGND 0.405233f
C756 VDPWR.n84 VGND 0.061913f
C757 VDPWR.n85 VGND 0.056913f
C758 VDPWR.n86 VGND 0.030855f
C759 VDPWR.n87 VGND 0.037021f
C760 VDPWR.n88 VGND 0.023938f
C761 VDPWR.n89 VGND 0.807609f
C762 VDPWR.t23 VGND 0.001565f
C763 VDPWR.t44 VGND 0.001565f
C764 VDPWR.n90 VGND 0.00313f
C765 VDPWR.n91 VGND 0.004476f
C766 VDPWR.t36 VGND 0.001565f
C767 VDPWR.t15 VGND 0.001565f
C768 VDPWR.n92 VGND 0.00313f
C769 VDPWR.n93 VGND 0.004476f
C770 VDPWR.n94 VGND 0.094814f
C771 VDPWR.t34 VGND 0.001565f
C772 VDPWR.t13 VGND 0.001565f
C773 VDPWR.n95 VGND 0.00313f
C774 VDPWR.n96 VGND 0.004476f
C775 VDPWR.t17 VGND 0.001565f
C776 VDPWR.t39 VGND 0.001565f
C777 VDPWR.n97 VGND 0.00313f
C778 VDPWR.n98 VGND 0.004476f
C779 VDPWR.n99 VGND 0.146582f
C780 VDPWR.t19 VGND 0.001565f
C781 VDPWR.t35 VGND 0.001565f
C782 VDPWR.n100 VGND 0.00313f
C783 VDPWR.n101 VGND 0.004476f
C784 VDPWR.t31 VGND 0.001565f
C785 VDPWR.t21 VGND 0.001565f
C786 VDPWR.n102 VGND 0.00313f
C787 VDPWR.n103 VGND 0.004476f
C788 VDPWR.n104 VGND 0.030697f
C789 VDPWR.n105 VGND 0.092284f
C790 VDPWR.t33 VGND 0.004533f
C791 VDPWR.t43 VGND 0.004533f
C792 VDPWR.n106 VGND 0.009293f
C793 VDPWR.n107 VGND 0.025644f
C794 VDPWR.n108 VGND 0.038921f
C795 VDPWR.n109 VGND 0.567005f
C796 VDPWR.n110 VGND 0.78771f
C797 VDPWR.n111 VGND 0.017906f
C798 VDPWR.n112 VGND 0.076846f
C799 VDPWR.n113 VGND 0.024591f
C800 VDPWR.n114 VGND 0.054924f
C801 VDPWR.n115 VGND 0.061618f
C802 VDPWR.n116 VGND 0.061618f
C803 VDPWR.n117 VGND 0.478933f
C804 VDPWR.t6 VGND 0.190001f
C805 VDPWR.t27 VGND 0.132715f
C806 VDPWR.t49 VGND 0.074358f
C807 VDPWR.t2 VGND 0.090359f
C808 VDPWR.t51 VGND 0.148716f
C809 VDPWR.t9 VGND 0.148716f
C810 VDPWR.t47 VGND 0.192013f
C811 VDPWR.t61 VGND 0.049545f
C812 VDPWR.t60 VGND 0.049545f
C813 VDPWR.n118 VGND 0.068002f
C814 VDPWR.n119 VGND 0.01319f
C815 VDPWR.n120 VGND 0.049068f
C816 VDPWR.n121 VGND 0.057729f
C817 VDPWR.n122 VGND 0.055525f
C818 VDPWR.n123 VGND 0.027565f
C819 VDPWR.n124 VGND 0.061913f
C820 VDPWR.n125 VGND 0.259805f
C821 VDPWR.n126 VGND 0.125237f
C822 VDPWR.t25 VGND 0.270154f
C823 VDPWR.t40 VGND 0.21587f
C824 VDPWR.n127 VGND 0.186521f
C825 VDPWR.t37 VGND 0.37276f
C826 VDPWR.n128 VGND 0.405233f
C827 VDPWR.n129 VGND 0.061913f
C828 VDPWR.n130 VGND 0.056913f
C829 VDPWR.n131 VGND 0.030855f
C830 VDPWR.n132 VGND 0.037021f
C831 flash_0.x7.pos_en_b.n0 VGND 0.766491f
C832 flash_0.x7.pos_en_b.t6 VGND 0.932199f
C833 flash_0.x7.pos_en_b.t4 VGND 0.216253f
C834 flash_0.x7.pos_en_b.t5 VGND 0.216253f
C835 flash_0.x7.pos_en_b.t3 VGND 0.010089f
C836 flash_0.x7.pos_en_b.t0 VGND 0.010089f
C837 flash_0.x7.pos_en_b.t1 VGND 0.008975f
C838 flash_0.x7.pos_en_b.n1 VGND 0.032452f
C839 flash_0.x7.pos_en_b.t2 VGND 0.008975f
C840 flash_0.x4.dcgint.t9 VGND 0.016015f
C841 flash_0.x4.dcgint.t10 VGND 0.016015f
C842 flash_0.x4.dcgint.t11 VGND 0.016015f
C843 flash_0.x4.dcgint.t5 VGND 0.017561f
C844 flash_0.x4.dcgint.n0 VGND 0.05401f
C845 flash_0.x4.dcgint.t3 VGND 0.017266f
C846 flash_0.x4.dcgint.t6 VGND 0.355987f
C847 flash_0.x4.dcgint.t0 VGND 0.222316f
C848 flash_0.x4.dcgint.t2 VGND 0.280884f
C849 flash_0.x4.dcgint.t1 VGND 0.004616f
C850 flash_0.x4.dcgint.t7 VGND 0.004616f
C851 flash_0.x4.dcgint.n1 VGND 0.009325f
C852 flash_0.x4.dcgint.t4 VGND 0.004616f
C853 flash_0.x4.dcgint.t8 VGND 0.004616f
C854 flash_0.x4.dcgint.n2 VGND 0.009325f
C855 flash_0.x4.dcgint.n3 VGND 0.045712f
C856 flash_0.x4.dcgint.n4 VGND 0.233815f
C857 flash_0.x4.dcgint.n5 VGND 0.046322f
C858 flash_0.x4.dcgint.n6 VGND 0.34091f
C859 flash_0.x4.VOUT.t8 VGND 0.00924f
C860 flash_0.x4.VOUT.t11 VGND 0.002436f
C861 flash_0.x4.VOUT.t10 VGND 0.002436f
C862 flash_0.x4.VOUT.n0 VGND 0.005005f
C863 flash_0.x4.VOUT.t13 VGND 0.002436f
C864 flash_0.x4.VOUT.t9 VGND 0.002436f
C865 flash_0.x4.VOUT.n1 VGND 0.005003f
C866 flash_0.x4.VOUT.t12 VGND 0.00924f
C867 flash_0.x4.VOUT.t7 VGND 0.008362f
C868 flash_0.x4.VOUT.t0 VGND 0.008358f
C869 flash_0.x4.VOUT.t14 VGND 0.099962f
C870 flash_0.x4.VOUT.t1 VGND 0.008626f
C871 flash_0.x4.VOUT.t4 VGND 0.008626f
C872 flash_0.x4.VOUT.t6 VGND 0.002436f
C873 flash_0.x4.VOUT.t3 VGND 0.002436f
C874 flash_0.x4.VOUT.n2 VGND 0.005003f
C875 flash_0.x4.VOUT.t2 VGND 0.002436f
C876 flash_0.x4.VOUT.t5 VGND 0.002436f
C877 flash_0.x4.VOUT.n3 VGND 0.005003f
C878 flash_0.x4.neg_mid_b.t10 VGND 0.828035f
C879 flash_0.x4.neg_mid_b.n0 VGND 0.140489f
C880 flash_0.x4.neg_mid_b.t2 VGND 0.027096f
C881 flash_0.x4.neg_mid_b.t4 VGND 0.007678f
C882 flash_0.x4.neg_mid_b.t5 VGND 0.007678f
C883 flash_0.x4.neg_mid_b.n1 VGND 0.015666f
C884 flash_0.x4.neg_mid_b.t9 VGND 0.085863f
C885 flash_0.x4.neg_mid_b.t6 VGND 0.02816f
C886 flash_0.x4.neg_mid_b.t3 VGND 0.02709f
C887 flash_0.x4.neg_mid_b.t7 VGND 0.067252f
C888 flash_0.x4.neg_mid_b.t8 VGND 0.122491f
C889 flash_0.x4.neg_mid_b.t12 VGND 0.067252f
C890 flash_0.x4.neg_mid_b.t14 VGND 0.122491f
C891 flash_0.x4.neg_mid_b.t11 VGND 0.067252f
C892 flash_0.x4.neg_mid_b.t13 VGND 0.122491f
C893 flash_0.x4.neg_mid_b.t1 VGND 0.007678f
C894 flash_0.x4.neg_mid_b.t0 VGND 0.007678f
C895 flash_0.x4.neg_mid_b.n2 VGND 0.015661f
C896 flash_0.x4.neg_en_b.n0 VGND 0.117521f
C897 flash_0.x4.neg_en_b.t2 VGND 0.036466f
C898 flash_0.x4.neg_en_b.t4 VGND 0.052338f
C899 flash_0.x4.neg_en_b.t8 VGND 0.051225f
C900 flash_0.x4.neg_en_b.t7 VGND 0.051225f
C901 flash_0.x4.neg_en_b.t5 VGND 0.051225f
C902 flash_0.x4.neg_en_b.t6 VGND 0.051201f
C903 flash_0.x4.neg_en_b.t9 VGND 0.051201f
C904 flash_0.x4.neg_en_b.t3 VGND 0.038945f
C905 flash_0.x4.neg_en_b.t0 VGND 0.032439f
C906 flash_0.x4.neg_en_b.t1 VGND 0.032439f
C907 ui_in[1].t17 VGND 0.038985f
C908 ui_in[1].n0 VGND 0.059558f
C909 ui_in[1].t10 VGND 0.038985f
C910 ui_in[1].n1 VGND 0.153802f
C911 ui_in[1].t12 VGND 0.038985f
C912 ui_in[1].n2 VGND 0.113223f
C913 ui_in[1].t13 VGND 0.038985f
C914 ui_in[1].n3 VGND 0.153802f
C915 ui_in[1].t15 VGND 0.038985f
C916 ui_in[1].n4 VGND 0.059558f
C917 ui_in[1].t2 VGND 0.038985f
C918 ui_in[1].n5 VGND 0.15152f
C919 ui_in[1].n6 VGND 0.421036f
C920 ui_in[1].t5 VGND 0.274588f
C921 ui_in[1].t0 VGND 0.286929f
C922 ui_in[1].n7 VGND 0.462789f
C923 ui_in[1].n8 VGND 0.341025f
C924 ui_in[1].t16 VGND 0.274588f
C925 ui_in[1].t14 VGND 0.286929f
C926 ui_in[1].n9 VGND 0.462789f
C927 ui_in[1].n10 VGND 0.234773f
C928 ui_in[1].n11 VGND 0.233332f
C929 ui_in[1].n12 VGND 0.131283f
C930 ui_in[1].n13 VGND 0.338374f
C931 ui_in[1].t7 VGND 0.229852f
C932 ui_in[1].t4 VGND 0.21134f
C933 ui_in[1].n14 VGND 0.323952f
C934 ui_in[1].n15 VGND 0.123876f
C935 ui_in[1].n16 VGND 0.167578f
C936 ui_in[1].t11 VGND 0.274588f
C937 ui_in[1].t8 VGND 0.286929f
C938 ui_in[1].n17 VGND 0.462789f
C939 ui_in[1].n18 VGND 0.230376f
C940 ui_in[1].n19 VGND 0.102431f
C941 ui_in[1].t9 VGND 0.274588f
C942 ui_in[1].t6 VGND 0.286929f
C943 ui_in[1].n20 VGND 0.462789f
C944 ui_in[1].n21 VGND 0.230376f
C945 ui_in[1].n22 VGND 0.103027f
C946 ui_in[1].n23 VGND 0.323672f
C947 ui_in[1].t3 VGND 0.229852f
C948 ui_in[1].t1 VGND 0.21134f
C949 ui_in[1].n24 VGND 0.323952f
C950 ui_in[1].n25 VGND 0.133376f
C951 ui_in[1].n26 VGND 0.524398f
C952 ui_in[1].n27 VGND 4.605279f
C953 ui_in[1].n28 VGND 0.525293f
C954 flash_0.x4.pos_mid_b.t0 VGND 0.019679f
C955 flash_0.x4.pos_mid_b.t1 VGND 0.019666f
C956 flash_0.x4.pos_mid_b.t8 VGND 0.055631f
C957 flash_0.x4.pos_mid_b.t7 VGND 0.055631f
C958 flash_0.x4.pos_mid_b.t4 VGND 0.055631f
C959 flash_0.x4.pos_mid_b.t3 VGND 0.055631f
C960 flash_0.x4.pos_mid_b.t6 VGND 0.055631f
C961 flash_0.x4.pos_mid_b.t5 VGND 0.055631f
C962 flash_0.x4.pos_mid_b.t2 VGND 0.020073f
C963 clk.t0 VGND 0.123904f
C964 clk.t1 VGND 0.116806f
C965 clk.n0 VGND 0.454326f
C966 clk.t2 VGND 0.123904f
C967 clk.t3 VGND 0.116806f
C968 clk.n1 VGND 0.454326f
C969 clk.n2 VGND 1.74152f
C970 clk.n3 VGND 4.1318f
C971 flash_0.x2.clkb.t0 VGND 0.011623f
C972 flash_0.x2.clkb.t1 VGND 0.018241f
C973 VAPWR.t14 VGND 0.003481f
C974 VAPWR.n0 VGND 0.025641f
C975 VAPWR.t1 VGND 0.003478f
C976 VAPWR.n1 VGND 0.034609f
C977 VAPWR.n2 VGND 0.04124f
C978 VAPWR.n3 VGND 0.025842f
C979 VAPWR.n4 VGND 0.045085f
C980 VAPWR.n5 VGND 0.148926f
C981 VAPWR.n6 VGND 0.050067f
C982 VAPWR.n7 VGND 0.050067f
C983 VAPWR.n8 VGND 0.022493f
C984 VAPWR.n9 VGND 0.022493f
C985 VAPWR.t15 VGND 0.010283f
C986 VAPWR.n10 VGND 0.022741f
C987 VAPWR.n11 VGND 0.130115f
C988 VAPWR.n12 VGND 0.130115f
C989 VAPWR.n13 VGND 0.183947f
C990 VAPWR.n14 VGND 0.049835f
C991 VAPWR.n15 VGND 0.022537f
C992 VAPWR.n16 VGND 0.030498f
C993 VAPWR.n17 VGND 0.022154f
C994 VAPWR.n18 VGND 0.020469f
C995 VAPWR.n19 VGND 0.030498f
C996 VAPWR.n20 VGND 0.022537f
C997 VAPWR.n21 VGND 0.048933f
C998 VAPWR.n22 VGND 0.030426f
C999 VAPWR.n23 VGND 0.022493f
C1000 VAPWR.n24 VGND 0.048933f
C1001 VAPWR.n25 VGND 0.190476f
C1002 VAPWR.n26 VGND 0.049075f
C1003 VAPWR.n27 VGND 0.183947f
C1004 VAPWR.n28 VGND 0.190476f
C1005 VAPWR.n29 VGND 0.183947f
C1006 VAPWR.n30 VGND 0.049075f
C1007 VAPWR.n31 VGND 0.016776f
C1008 VAPWR.n32 VGND 0.016833f
C1009 VAPWR.n33 VGND 0.022071f
C1010 VAPWR.n34 VGND 0.147307f
C1011 VAPWR.n35 VGND 0.020469f
C1012 VAPWR.n36 VGND 0.030498f
C1013 VAPWR.n37 VGND 0.022537f
C1014 VAPWR.n38 VGND 0.048933f
C1015 VAPWR.n39 VGND 0.030426f
C1016 VAPWR.n40 VGND 0.022493f
C1017 VAPWR.n41 VGND 0.049459f
C1018 VAPWR.n42 VGND 0.190476f
C1019 VAPWR.n43 VGND 0.049143f
C1020 VAPWR.n44 VGND 0.183947f
C1021 VAPWR.n45 VGND 0.190476f
C1022 VAPWR.n46 VGND 0.183947f
C1023 VAPWR.n47 VGND 0.049143f
C1024 VAPWR.n48 VGND 0.016776f
C1025 VAPWR.n49 VGND 0.016833f
C1026 VAPWR.n50 VGND 0.022071f
C1027 VAPWR.n51 VGND 0.034828f
C1028 VAPWR.n52 VGND 0.306925f
C1029 VAPWR.n53 VGND 0.083428f
C1030 VAPWR.n54 VGND 0.054859f
C1031 VAPWR.n55 VGND 0.073402f
C1032 VAPWR.n56 VGND 0.028091f
C1033 VAPWR.n57 VGND 0.022537f
C1034 VAPWR.n58 VGND 0.049832f
C1035 VAPWR.n59 VGND 0.15277f
C1036 VAPWR.n60 VGND 0.188825f
C1037 VAPWR.n61 VGND 0.135464f
C1038 VAPWR.n62 VGND 0.033985f
C1039 VAPWR.n63 VGND 0.015983f
C1040 VAPWR.t2 VGND 0.037542f
C1041 VAPWR.t13 VGND 0.343435f
C1042 VAPWR.t0 VGND 0.182547f
C1043 VAPWR.n64 VGND 0.142205f
C1044 VAPWR.n65 VGND 0.019665f
C1045 VAPWR.n66 VGND 0.026555f
C1046 VAPWR.n67 VGND 0.00647f
C1047 VAPWR.t3 VGND 0.010229f
C1048 VAPWR.n68 VGND 0.055175f
C1049 VAPWR.n69 VGND 0.059815f
C1050 VAPWR.n70 VGND 0.096071f
C1051 VAPWR.t12 VGND 0.003478f
C1052 VAPWR.n71 VGND 0.017733f
C1053 VAPWR.t5 VGND 0.003481f
C1054 VAPWR.n72 VGND 0.025711f
C1055 VAPWR.n73 VGND 0.045085f
C1056 VAPWR.n74 VGND 0.148926f
C1057 VAPWR.n75 VGND 0.050067f
C1058 VAPWR.n76 VGND 0.050067f
C1059 VAPWR.n77 VGND 0.022493f
C1060 VAPWR.n78 VGND 0.022493f
C1061 VAPWR.t7 VGND 0.010283f
C1062 VAPWR.n79 VGND 0.121994f
C1063 VAPWR.n80 VGND 0.01091f
C1064 VAPWR.n81 VGND 0.018798f
C1065 VAPWR.n82 VGND 0.011001f
C1066 VAPWR.n83 VGND 0.018798f
C1067 VAPWR.n84 VGND 0.085518f
C1068 VAPWR.t9 VGND 0.104521f
C1069 VAPWR.n87 VGND 0.085518f
C1070 VAPWR.t10 VGND 0.006509f
C1071 VAPWR.n88 VGND 0.040216f
C1072 VAPWR.n89 VGND 0.13191f
C1073 VAPWR.n90 VGND 0.065256f
C1074 VAPWR.n91 VGND 0.130115f
C1075 VAPWR.n92 VGND 0.130115f
C1076 VAPWR.n93 VGND 0.183947f
C1077 VAPWR.n94 VGND 0.049835f
C1078 VAPWR.n95 VGND 0.023894f
C1079 VAPWR.n96 VGND 0.094738f
C1080 VAPWR.t8 VGND 0.019586f
C1081 VAPWR.n97 VGND 0.006748f
C1082 VAPWR.n98 VGND 0.003219f
C1083 VAPWR.n99 VGND 0.057898f
C1084 VAPWR.n100 VGND 0.081102f
C1085 VAPWR.n101 VGND 0.023469f
C1086 VAPWR.n102 VGND 0.038288f
C1087 VAPWR.n103 VGND 0.030914f
C1088 VAPWR.n104 VGND 0.005625f
C1089 VAPWR.n105 VGND 0.027268f
C1090 VAPWR.n106 VGND 0.01091f
C1091 VAPWR.n107 VGND 0.011001f
C1092 VAPWR.n108 VGND 0.018067f
C1093 VAPWR.n109 VGND 0.022537f
C1094 VAPWR.n110 VGND 0.049832f
C1095 VAPWR.n111 VGND 0.15277f
C1096 VAPWR.n112 VGND 0.188825f
C1097 VAPWR.n113 VGND 0.135464f
C1098 VAPWR.n114 VGND 0.033985f
C1099 VAPWR.n115 VGND 0.015983f
C1100 VAPWR.t6 VGND 0.037542f
C1101 VAPWR.t4 VGND 0.343435f
C1102 VAPWR.t11 VGND 0.182547f
C1103 VAPWR.n116 VGND 0.142205f
C1104 VAPWR.n117 VGND 0.019665f
C1105 VAPWR.n118 VGND 0.026555f
C1106 VAPWR.n119 VGND 0.018775f
C1107 VAPWR.t16 VGND 0.010259f
C1108 VAPWR.n120 VGND 0.094854f
C1109 VAPWR.n121 VGND 0.11419f
C1110 VAPWR.n122 VGND 0.018245f
C1111 VAPWR.n123 VGND 1.0575f
C1112 VAPWR.n124 VGND 0.521869f
C1113 VAPWR.n125 VGND 7.2806f
C1114 VAPWR.n126 VGND 40.983803f
C1115 flash_0.x7.VPRGPOS.t26 VGND 0.001628f
C1116 flash_0.x7.VPRGPOS.t20 VGND 0.048001f
C1117 flash_0.x7.VPRGPOS.t13 VGND 0.030458f
C1118 flash_0.x7.VPRGPOS.t14 VGND 0.030458f
C1119 flash_0.x7.VPRGPOS.t18 VGND 0.030458f
C1120 flash_0.x7.VPRGPOS.t15 VGND 0.02988f
C1121 flash_0.x7.VPRGPOS.t22 VGND 0.130893f
C1122 flash_0.x7.VPRGPOS.t16 VGND 0.050507f
C1123 flash_0.x7.VPRGPOS.n0 VGND 0.006722f
C1124 flash_0.x7.VPRGPOS.t23 VGND 0.001628f
C1125 flash_0.x7.VPRGPOS.t30 VGND 0.001628f
C1126 flash_0.x7.VPRGPOS.t10 VGND 0.003253f
C1127 flash_0.x7.VPRGPOS.t9 VGND 0.001739f
C1128 flash_0.x7.VPRGPOS.n1 VGND 0.025524f
C1129 flash_0.x7.VPRGPOS.n2 VGND 0.025599f
C1130 flash_0.x7.VPRGPOS.n4 VGND 0.043977f
C1131 flash_0.x7.VPRGPOS.n5 VGND 0.026181f
C1132 flash_0.x7.VPRGPOS.n6 VGND 0.300528f
C1133 flash_0.x7.VPRGPOS.t8 VGND 0.482339f
C1134 flash_0.x7.VPRGPOS.n8 VGND 0.043977f
C1135 flash_0.x7.VPRGPOS.n9 VGND 0.300528f
C1136 flash_0.x7.VPRGPOS.n10 VGND 0.014456f
C1137 flash_0.x7.VPRGPOS.n11 VGND 0.014476f
C1138 flash_0.x7.VPRGPOS.n12 VGND 0.030642f
C1139 flash_0.x7.VPRGPOS.t32 VGND 0.001628f
C1140 flash_0.x7.VPRGPOS.t7 VGND 4.6e-19
C1141 flash_0.x7.VPRGPOS.t3 VGND 4.6e-19
C1142 flash_0.x7.VPRGPOS.n13 VGND 9.44e-19
C1143 flash_0.x7.VPRGPOS.t12 VGND 4.6e-19
C1144 flash_0.x7.VPRGPOS.t1 VGND 4.6e-19
C1145 flash_0.x7.VPRGPOS.n14 VGND 9.44e-19
C1146 flash_0.x7.VPRGPOS.t31 VGND 0.001628f
C1147 flash_0.x7.VPRGPOS.t17 VGND 0.048001f
C1148 flash_0.x7.VPRGPOS.t6 VGND 0.030458f
C1149 flash_0.x7.VPRGPOS.t2 VGND 0.030458f
C1150 flash_0.x7.VPRGPOS.t11 VGND 0.030458f
C1151 flash_0.x7.VPRGPOS.t0 VGND 0.02988f
C1152 flash_0.x7.VPRGPOS.t4 VGND 0.130893f
C1153 flash_0.x7.VPRGPOS.t19 VGND 0.050507f
C1154 flash_0.x7.VPRGPOS.n15 VGND 0.006722f
C1155 flash_0.x7.VPRGPOS.t5 VGND 0.001628f
C1156 flash_0.x7.VPRGPOS.t29 VGND 0.001628f
C1157 flash_0.x7.VPRGPOS.n16 VGND 0.115389f
C1158 flash_0.x7.VPRGPOS.n17 VGND 1.98663f
C1159 flash_0.x7.VPRGPOS.t24 VGND 0.001628f
C1160 flash_0.x7.VPRGPOS.t25 VGND 4.6e-19
C1161 flash_0.x7.VPRGPOS.t21 VGND 4.6e-19
C1162 flash_0.x7.VPRGPOS.n18 VGND 9.44e-19
C1163 flash_0.x7.VPRGPOS.t27 VGND 4.6e-19
C1164 flash_0.x7.VPRGPOS.t28 VGND 4.6e-19
C1165 flash_0.x7.VPRGPOS.n19 VGND 9.44e-19
C1166 flash_0.x7.pos_mid_b.t0 VGND 0.020534f
C1167 flash_0.x7.pos_mid_b.t1 VGND 0.020521f
C1168 flash_0.x7.pos_mid_b.t5 VGND 0.05805f
C1169 flash_0.x7.pos_mid_b.t4 VGND 0.05805f
C1170 flash_0.x7.pos_mid_b.t3 VGND 0.05805f
C1171 flash_0.x7.pos_mid_b.t6 VGND 0.05805f
C1172 flash_0.x7.pos_mid_b.t8 VGND 0.05805f
C1173 flash_0.x7.pos_mid_b.t7 VGND 0.05805f
C1174 flash_0.x7.pos_mid_b.t2 VGND 0.020946f
.ends

