* NGSPICE file created from flash.ext - technology: sky130A

.subckt charge_pump VAPWR VOUT clk VGND stage2 stage1
X0 clkina clkinb VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X1 clkinb clk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X2 stage1 VAPWR VAPWR VAPWR sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 stage2 stage1 stage1 stage1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 clkb clkinb VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X5 clkb clkinb VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X6 VOUT VGND sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X7 VOUT stage2 stage2 stage2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X8 clkinb clk VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X9 clkina clkinb VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X10 clka clkina VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X11 clkb stage2 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X12 clka clkina VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X13 clka stage1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
.ends

.subckt charge_pump_neg_nmos clk VOUT VAPWR VGND stage2 stage1
X0 clkina clkinb VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X1 clkinb clk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X2 stage1 stage1 VGND stage1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 stage2 stage2 stage1 stage2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 clkb clkinb VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X5 clkb clkinb VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X6 VOUT VGND sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X7 VOUT VOUT stage2 VOUT sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X8 clkinb clk VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X9 clkina clkinb VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X10 clka clkina VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X11 clkb stage2 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X12 clka clkina VAPWR VAPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X13 clka stage1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
.ends

.subckt vprog_controller pos_en neg_en VOUT VGND VPRGPOS VPRGNEG VDPWR VDPWR1
X0 VDPWR neg_en neg_mid VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X1 pos_mid_b pos_en VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X2 VOUT neg_mid_b dcgint dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X3 VDPWR pos_en pos_en_b VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X4 VOUT VDPWR1 vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X5 dcgint neg_mid_b VOUT dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X6 pos_mid_b pos_en VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X7 vintp pos_mid_b VPRGPOS VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X8 neg_en_b neg_en VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X9 VPRGPOS pos_mid_b vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X10 VOUT neg_mid_b dcgint dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X11 dcgint neg_mid_b VOUT dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X12 pos_mid pos_en_b VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X13 neg_en_b neg_en VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=3
X14 neg_mid neg_en VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X15 vintp pos_mid_b VPRGPOS VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X16 VDPWR neg_en_b neg_mid_b VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X17 VDPWR neg_en_b neg_mid_b VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X18 a_2408_n3852# neg_mid_b VPRGNEG VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X19 VDPWR neg_en_b neg_mid_b VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X20 neg_mid neg_en VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X21 vintp VDPWR1 VOUT VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X22 pos_mid pos_en_b VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X23 neg_mid neg_en VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X24 VOUT VDPWR1 vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X25 VGND pos_en_b pos_mid VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X26 pos_en_b pos_en VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X27 a_2408_n3852# neg_mid_b VPRGNEG VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X28 vintp VDPWR1 VOUT VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X29 VGND pos_en_b pos_mid VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X30 pos_en_b pos_en VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X31 VPRGPOS pos_mid_b vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X32 VGND neg_en neg_en_b VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X33 vintp pos_mid_b VPRGPOS VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X34 dcgint pos_en_b VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X35 VDPWR neg_en neg_mid VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X36 VDPWR neg_en neg_en_b VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X37 VDPWR neg_en neg_mid VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X38 dcgint pos_en_b VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X39 VPRGPOS pos_mid pos_mid_b VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X40 neg_mid_b neg_mid VPRGNEG VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=1
X41 neg_mid_b neg_en_b VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X42 neg_mid_b neg_en_b VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X43 VOUT VDPWR1 vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X44 VPRGNEG neg_mid_b neg_mid VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.145 ps=1.58 w=0.5 l=1
X45 dcgint neg_mid_b VOUT dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X46 vintp VDPWR1 VOUT VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X47 VGND pos_en pos_mid_b VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X48 VOUT VDPWR a_2408_n3852# VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X49 dcgint pos_en_b VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X50 VPRGPOS pos_mid_b pos_mid VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X51 VGND pos_en pos_mid_b VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X52 VOUT VDPWR a_2408_n3852# VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X53 VPRGPOS pos_mid_b vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X54 neg_mid_b neg_en_b VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X55 dcgint neg_mid_b VOUT dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X56 VGND pos_en pos_en_b VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
.ends

.subckt sky130_fd_pr__pfet_01v8_29FY9H a_n300_n197# a_300_n100# a_n358_n100# w_n496_n319#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n496_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__nfet_01v8_KAAY2V a_300_n100# a_n358_n100# a_n300_n188# a_n460_n274#
X0 a_300_n100# a_n300_n188# a_n358_n100# a_n460_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt inverter A Y VDD VSS
XXM1 A Y VDD VDD sky130_fd_pr__pfet_01v8_29FY9H
XXM2 Y VSS A VSS sky130_fd_pr__nfet_01v8_KAAY2V
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_VPAE37 a_n2058_n50# a_n2000_n147# a_2000_n50#
+ w_n2258_n347#
X0 a_2000_n50# a_n2000_n147# a_n2058_n50# w_n2258_n347# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_GJ3XY6 a_1000_n50# w_n1258_n347# a_n1000_n147#
+ a_n1058_n50#
X0 a_1000_n50# a_n1000_n147# a_n1058_n50# w_n1258_n347# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=10
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_9UU773 a_50_n500# a_n242_n722# a_n108_n500# a_n50_n588#
X0 a_50_n500# a_n50_n588# a_n108_n500# a_n242_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_HQS8YU a_50_n200# a_n242_n422# a_n108_n200# a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_bs_flash__special_sonosfet_star_EA7MKQ a_n83_n45# dw_n439_n473#
+ a_n33_n133# a_22_n45# w_n439_n473#
X0 a_22_n45# a_n33_n133# a_n83_n45# w_n439_n473# sky130_fd_bs_flash__special_sonosfet_star ad=0.13725 pd=1.51 as=0.13725 ps=1.51 w=0.45 l=0.22
.ends

.subckt flash VDPWR VAPWR VGND clk prog_en erase_en read_en data_out VPROGMON
Xx3 VAPWR x3/VOUT clk VGND x3/stage2 x3/stage1 charge_pump
Xx2 clk x2/VOUT VAPWR VGND x2/stage2 x2/stage1 charge_pump_neg_nmos
Xx4 prog_en erase_en x4/VOUT VGND x3/VOUT x2/VOUT VDPWR VDPWR vprog_controller
Xx5 x5/A data_out VDPWR VGND inverter
Xx6 read_en x6/Y VDPWR VGND inverter
Xx7 erase_en prog_en x7/VOUT VGND x3/VOUT x2/VOUT VDPWR VDPWR vprog_controller
XXM1 li_7306_n1074# li_7306_n1074# x3/VOUT x3/VOUT sky130_fd_pr__pfet_g5v0d10v5_VPAE37
XXM2 VPROGMON VPROGMON li_7306_n1074# li_7306_n1074# sky130_fd_pr__pfet_g5v0d10v5_VPAE37
XXM3 VPROGMON VPROGMON VGND VGND sky130_fd_pr__pfet_g5v0d10v5_GJ3XY6
XXM4 VDPWR x6/Y x5/A VDPWR sky130_fd_pr__pfet_g5v0d10v5_VPAE37
XXM5 x5/A x5/A m1_4558_2458# x5/A sky130_fd_pr__nfet_g5v0d10v5_9UU773
XXM8 m1_2666_2466# VGND VGND read_en sky130_fd_pr__nfet_g5v0d10v5_HQS8YU
XX1 m1_2666_2466# x3/VOUT x4/VOUT m1_4558_2458# x7/VOUT sky130_fd_bs_flash__special_sonosfet_star_EA7MKQ
.ends

