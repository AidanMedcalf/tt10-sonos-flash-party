magic
tech sky130A
magscale 1 2
timestamp 1740014482
<< error_s >>
rect 10490 2670 10548 2676
rect 10490 2636 10502 2670
rect 10490 2630 10548 2636
rect 10497 2508 10541 2598
rect 10490 2470 10548 2476
rect 10490 2436 10502 2470
rect 10490 2430 10548 2436
<< nwell >>
rect 9800 2816 11238 3306
rect 9800 2290 10290 2816
rect 10748 2290 11238 2816
rect 9800 1800 11238 2290
<< mvnsubdiff >>
rect 10000 2064 10088 2088
rect 10000 2024 10024 2064
rect 10064 2024 10088 2064
rect 10000 2000 10088 2024
<< mvnsubdiffcont >>
rect 10024 2024 10064 2064
<< locali >>
rect 10008 2064 10080 2080
rect 10008 2024 10024 2064
rect 10064 2024 10080 2064
rect 10008 2008 10080 2024
use sky130_fd_bs_flash__special_sonosfet_star_EA7MKQ  X1
timestamp 1739996772
transform 1 0 10519 0 1 2553
box -519 -553 519 553
use charge_pump_neg_nmos  x2 ../charge_pump_neg_nmos
timestamp 1739484054
transform 1 0 4288 0 1 11688
box -4288 -1488 12990 4458
use charge_pump  x3 ../charge_pump
timestamp 1739252499
transform 1 0 4288 0 1 5488
box -4288 -1488 12990 4458
use vprog_controller  x4 ../vprog_controller
timestamp 1738900598
transform 1 0 14676 0 1 10282
box 1324 -4282 4846 -1260
use inverter  x5 ../inverter
timestamp 1739087840
transform 1 0 16000 0 1 2620
box 0 -620 992 638
use inverter  x6
timestamp 1739087840
transform 1 0 0 0 1 2620
box 0 -620 992 638
use vprog_controller  x7
timestamp 1738900598
transform 1 0 14676 0 1 16282
box 1324 -4282 4846 -1260
use sky130_fd_pr__pfet_g5v0d10v5_VPAE37  XM1
timestamp 1739996415
transform 1 0 2258 0 1 347
box -2258 -347 2258 347
use sky130_fd_pr__pfet_g5v0d10v5_VPAE37  XM2
timestamp 1739996415
transform 1 0 6774 0 1 347
box -2258 -347 2258 347
use sky130_fd_pr__pfet_g5v0d10v5_GJ3XY6  XM3
timestamp 1739996415
transform 1 0 10290 0 1 347
box -1258 -347 1258 347
use sky130_fd_pr__pfet_g5v0d10v5_VPAE37  XM4
timestamp 1739996415
transform 1 0 4258 0 1 2347
box -2258 -347 2258 347
use sky130_fd_pr__nfet_g5v0d10v5_9UU773  XM5
timestamp 1739996415
transform 1 0 8278 0 1 2758
box -278 -758 278 758
use sky130_fd_pr__nfet_g5v0d10v5_HQS8YU  XM8
timestamp 1739996415
transform 1 0 14278 0 1 2458
box -278 -458 278 458
<< end >>
