magic
tech sky130A
magscale 1 2
timestamp 1739996415
<< nwell >>
rect -2258 -347 2258 347
<< mvpmos >>
rect -2000 -50 2000 50
<< mvpdiff >>
rect -2058 38 -2000 50
rect -2058 -38 -2046 38
rect -2012 -38 -2000 38
rect -2058 -50 -2000 -38
rect 2000 38 2058 50
rect 2000 -38 2012 38
rect 2046 -38 2058 38
rect 2000 -50 2058 -38
<< mvpdiffc >>
rect -2046 -38 -2012 38
rect 2012 -38 2046 38
<< mvnsubdiff >>
rect -2192 269 2192 281
rect -2192 235 -2084 269
rect 2084 235 2192 269
rect -2192 223 2192 235
rect -2192 173 -2134 223
rect -2192 -173 -2180 173
rect -2146 -173 -2134 173
rect 2134 173 2192 223
rect -2192 -223 -2134 -173
rect 2134 -173 2146 173
rect 2180 -173 2192 173
rect 2134 -223 2192 -173
rect -2192 -235 2192 -223
rect -2192 -269 -2084 -235
rect 2084 -269 2192 -235
rect -2192 -281 2192 -269
<< mvnsubdiffcont >>
rect -2084 235 2084 269
rect -2180 -173 -2146 173
rect 2146 -173 2180 173
rect -2084 -269 2084 -235
<< poly >>
rect -2000 131 2000 147
rect -2000 97 -1984 131
rect 1984 97 2000 131
rect -2000 50 2000 97
rect -2000 -97 2000 -50
rect -2000 -131 -1984 -97
rect 1984 -131 2000 -97
rect -2000 -147 2000 -131
<< polycont >>
rect -1984 97 1984 131
rect -1984 -131 1984 -97
<< locali >>
rect -2180 235 -2084 269
rect 2084 235 2180 269
rect -2180 173 -2146 235
rect 2146 173 2180 235
rect -2000 97 -1984 131
rect 1984 97 2000 131
rect -2046 38 -2012 54
rect -2046 -54 -2012 -38
rect 2012 38 2046 54
rect 2012 -54 2046 -38
rect -2000 -131 -1984 -97
rect 1984 -131 2000 -97
rect -2180 -235 -2146 -173
rect 2146 -235 2180 -173
rect -2180 -269 -2084 -235
rect 2084 -269 2180 -235
<< viali >>
rect -1984 97 1984 131
rect -2046 -38 -2012 38
rect 2012 -38 2046 38
rect -1984 -131 1984 -97
<< metal1 >>
rect -1996 131 1996 137
rect -1996 97 -1984 131
rect 1984 97 1996 131
rect -1996 91 1996 97
rect -2052 38 -2006 50
rect -2052 -38 -2046 38
rect -2012 -38 -2006 38
rect -2052 -50 -2006 -38
rect 2006 38 2052 50
rect 2006 -38 2012 38
rect 2046 -38 2052 38
rect 2006 -50 2052 -38
rect -1996 -97 1996 -91
rect -1996 -131 -1984 -97
rect 1984 -131 1996 -97
rect -1996 -137 1996 -131
<< properties >>
string FIXED_BBOX -2163 -252 2163 252
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 20.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 ad {int((nf+1)/2) * W/nf * 0.29} as {int((nf+2)/2) * W/nf * 0.29} pd {2*int((nf+1)/2) * (W/nf + 0.29)} ps {2*int((nf+2)/2) * (W/nf + 0.29)} nrd {0.29 / W} nrs {0.29 / W} sa 0 sb 0 sd 0 mult 1
<< end >>
