magic
tech sky130A
magscale 1 2
timestamp 1740650923
<< error_s >>
rect 4496 2437 4540 2527
<< dnwell >>
rect 6050 3038 7044 3462
rect 6048 2962 7044 3038
rect 4756 2002 7044 2962
rect 6034 1928 7044 2002
rect 6050 1512 7044 1928
<< nwell >>
rect 5789 3242 7125 3542
rect 5789 3235 6280 3242
rect 3799 2745 6280 3235
rect 3799 2219 4289 2745
rect 4747 2219 6280 2745
rect 3799 1752 6280 2219
rect 5904 1726 6280 1752
rect 6836 3031 7125 3242
rect 6836 1726 7124 3031
rect 5904 1362 7124 1726
<< mvnsubdiff >>
rect 4974 3124 5116 3148
rect 4974 3038 4998 3124
rect 5092 3038 5116 3124
rect 4974 3014 5116 3038
<< mvnsubdiffcont >>
rect 4998 3038 5092 3124
<< locali >>
rect 4974 3138 5116 3148
rect 4974 3038 4990 3138
rect 5104 3038 5116 3138
rect 4974 3014 5116 3038
<< viali >>
rect 4990 3124 5104 3138
rect 4990 3038 4998 3124
rect 4998 3038 5092 3124
rect 5092 3038 5104 3124
rect 2368 2540 2406 2858
rect 4416 2668 4612 2706
rect 4330 2568 4364 2638
rect 4670 2568 4704 2638
rect 6746 1874 6786 3092
rect 4380 44 4430 406
rect 2390 -1058 2448 -674
rect 7306 -1074 7360 -672
rect 12228 -1046 12280 -678
<< metal1 >>
rect 12144 13506 12154 13518
rect 11706 13364 12154 13506
rect 12412 13506 12422 13518
rect 14248 13506 14392 13510
rect 12412 13364 14392 13506
rect 11706 13362 14392 13364
rect 3450 12528 5382 12728
rect 3450 9990 3650 12528
rect 3748 12027 3848 12042
rect 3748 11927 5284 12027
rect 3438 9984 3662 9990
rect 3438 9784 3450 9984
rect 3650 9784 3662 9984
rect 3438 9778 3662 9784
rect 3748 7690 3848 11927
rect 3931 9771 3941 9981
rect 4151 9771 5390 9981
rect 112 7590 122 7690
rect 222 7590 3848 7690
rect 3748 5998 3848 7590
rect 5180 6492 5390 9771
rect 3748 5898 5286 5998
rect 14248 4038 14392 13362
rect 4976 3894 14392 4038
rect 2340 3168 2350 3260
rect 2442 3168 2452 3260
rect 2350 2858 2442 3168
rect 4976 3138 5120 3894
rect 4976 3038 4990 3138
rect 5104 3038 5120 3138
rect 4976 3014 5120 3038
rect 6136 3428 14110 3508
rect 2350 2540 2368 2858
rect 2406 2600 2442 2858
rect 2406 2540 2534 2600
rect 2350 2508 2534 2540
rect 2581 2298 2609 2801
rect 4310 2706 4730 2734
rect 4310 2668 4416 2706
rect 4612 2668 4730 2706
rect 4310 2654 4730 2668
rect 4310 2638 4390 2654
rect 4310 2568 4330 2638
rect 4364 2568 4390 2638
rect 4650 2638 4730 2654
rect 4462 2568 4472 2622
rect 4538 2568 4548 2622
rect 4650 2568 4670 2638
rect 4704 2634 4730 2638
rect 6136 2634 6216 3428
rect 6740 3092 6792 3104
rect 6532 3026 6672 3058
rect 4704 2568 6216 2634
rect 4310 2558 4390 2568
rect 4324 2556 4370 2558
rect 4650 2554 6216 2568
rect 2666 2466 4466 2502
rect 4558 2458 6478 2498
rect 4460 2344 4470 2400
rect 4544 2344 4554 2400
rect 6640 2392 6672 3026
rect 6740 2392 6746 3092
rect 6640 2334 6746 2392
rect 2562 2072 2626 2298
rect 14 2010 2626 2072
rect 14 2008 2622 2010
rect 14 1214 78 2008
rect 6640 1946 6672 2334
rect 424 1826 2044 1946
rect 6568 1914 6672 1946
rect 6740 1874 6746 2334
rect 6786 2392 6792 3092
rect 7468 2624 7478 2718
rect 7572 2716 7582 2718
rect 7572 2624 8138 2716
rect 6786 2334 8483 2392
rect 6786 1874 6792 2334
rect 6740 1862 6792 1874
rect 6746 1834 6792 1862
rect 424 1790 544 1826
rect 116 1670 126 1790
rect 246 1670 578 1790
rect 458 1550 578 1670
rect 458 1430 1041 1550
rect 1924 1406 2044 1826
rect 1924 1286 4068 1406
rect 14 1150 274 1214
rect 338 1150 1379 1214
rect 1690 1150 3904 1214
rect 682 896 1032 900
rect 682 844 692 896
rect 744 844 1032 896
rect 682 836 1032 844
rect 756 -848 820 836
rect 3840 -270 3904 1150
rect 3948 290 4068 1286
rect 7261 1259 7319 2334
rect 8792 2330 8992 2394
rect 9056 2330 9066 2394
rect 7980 2018 7990 2080
rect 8136 2018 8146 2080
rect 7261 1201 8895 1259
rect 7261 1191 7319 1201
rect 4374 406 4436 418
rect 4374 290 4380 406
rect 3948 170 4380 290
rect 4374 44 4380 170
rect 4430 290 4436 406
rect 4430 170 4554 290
rect 4430 44 4436 170
rect 4374 32 4436 44
rect 5048 -270 5112 364
rect 8837 247 8895 1201
rect 14030 996 14110 3428
rect 14020 916 14030 996
rect 14110 916 14120 996
rect 12758 712 12768 764
rect 12832 712 12842 764
rect 12778 448 12820 712
rect 12778 412 13720 448
rect 14248 346 14392 3894
rect 16878 710 16888 762
rect 16952 710 16962 762
rect 16904 444 16946 710
rect 16904 412 17844 444
rect 8569 189 8895 247
rect 11236 202 11246 346
rect 11390 202 15364 346
rect 8837 169 8895 189
rect 3840 -334 5112 -270
rect 2384 -674 2456 -584
rect 2384 -828 2390 -674
rect 190 -912 820 -848
rect 2274 -912 2390 -828
rect 756 -1046 820 -912
rect 2384 -1058 2390 -912
rect 2448 -828 2456 -674
rect 7294 -672 7372 -622
rect 3120 -828 3282 -710
rect 7294 -822 7306 -672
rect 2448 -834 3282 -828
rect 2448 -904 2526 -834
rect 2856 -904 3282 -834
rect 2448 -912 3282 -904
rect 2448 -1058 2456 -912
rect 3120 -1024 3282 -912
rect 7166 -920 7306 -822
rect 2384 -1160 2456 -1058
rect 7294 -1074 7306 -920
rect 7360 -822 7372 -672
rect 12216 -678 12294 -654
rect 8026 -822 8178 -704
rect 12216 -820 12228 -678
rect 7360 -920 8178 -822
rect 7360 -1074 7372 -920
rect 8026 -1036 8178 -920
rect 12088 -922 12228 -820
rect 12216 -1046 12228 -922
rect 12280 -820 12294 -678
rect 12647 -820 12749 202
rect 15354 200 15364 202
rect 15506 202 15520 346
rect 15506 200 15516 202
rect 12280 -922 12749 -820
rect 12280 -1046 12294 -922
rect 12216 -1056 12294 -1046
rect 12222 -1058 12286 -1056
rect 7294 -1112 7372 -1074
<< via1 >>
rect 12154 13364 12412 13518
rect 3450 9784 3650 9984
rect 3941 9771 4151 9981
rect 122 7590 222 7690
rect 2350 3168 2442 3260
rect 4472 2568 4538 2622
rect 4470 2344 4544 2400
rect 7478 2624 7572 2718
rect 126 1670 246 1790
rect 274 1150 338 1214
rect 692 844 744 896
rect 8992 2330 9056 2394
rect 7990 2018 8136 2080
rect 14030 916 14110 996
rect 12768 712 12832 764
rect 16888 710 16952 762
rect 11246 202 11390 346
rect 2526 -904 2856 -834
rect 15364 200 15506 346
<< metal2 >>
rect 11520 13518 12412 13542
rect 11520 13366 12154 13518
rect 12154 13354 12412 13364
rect 4802 11341 5572 11541
rect -103 9991 4114 10040
rect -103 9984 4151 9991
rect -103 9784 3450 9984
rect 3650 9981 4151 9984
rect 3650 9784 3941 9981
rect -103 9771 3941 9784
rect -103 9761 4151 9771
rect -103 9640 4114 9761
rect -75 7690 325 7764
rect -75 7590 122 7690
rect 222 7590 325 7690
rect -75 7364 325 7590
rect 4802 5512 5002 11341
rect 11536 7342 11929 7528
rect 4802 5312 5650 5512
rect -12 3464 3608 3496
rect 4802 3464 5002 5312
rect 11743 3733 11929 7342
rect 10679 3547 14957 3733
rect -12 3264 10306 3464
rect -12 3260 3608 3264
rect -12 3168 2350 3260
rect 2442 3168 3608 3260
rect -12 3096 3608 3168
rect -37 1878 363 1929
rect -37 1868 606 1878
rect -37 1790 350 1868
rect -37 1670 126 1790
rect 246 1670 350 1790
rect -37 1612 350 1670
rect -37 1602 606 1612
rect -37 1529 363 1602
rect -22 1214 378 1333
rect -22 1150 274 1214
rect 338 1150 378 1214
rect -22 933 378 1150
rect 680 896 754 3096
rect 7478 2718 7572 2728
rect 4464 2632 4536 2634
rect 4464 2622 4538 2632
rect 4464 2568 4472 2622
rect 4464 2558 4538 2568
rect 4464 2410 4536 2558
rect 4464 2400 4544 2410
rect 4464 2344 4470 2400
rect 4464 2334 4544 2344
rect 4464 1524 4536 2334
rect 7478 1804 7572 2624
rect 7662 2086 7728 3264
rect 8974 2394 9374 2584
rect 8974 2330 8992 2394
rect 9056 2330 9374 2394
rect 8974 2184 9374 2330
rect 10106 2568 10306 3264
rect 10679 2739 10865 3547
rect 11004 3290 14252 3490
rect 11004 2568 11204 3290
rect 14052 3144 14252 3290
rect 13564 2944 14252 3144
rect 10106 2368 11204 2568
rect 14052 2506 14252 2944
rect 14771 2733 14957 3547
rect 15160 3550 17898 3750
rect 15160 2506 15360 3550
rect 17698 2954 17898 3550
rect 7990 2086 8136 2090
rect 7662 2080 8141 2086
rect 7662 2020 7990 2080
rect 8136 2020 8141 2080
rect 7990 2008 8136 2018
rect 7478 1694 7572 1704
rect 4464 1452 9326 1524
rect 680 844 692 896
rect 744 844 754 896
rect 680 834 754 844
rect 9254 186 9326 1452
rect 10106 1410 10306 2368
rect 14052 2306 15360 2506
rect 11218 1930 11418 1940
rect 11218 1792 11418 1802
rect 12752 1930 12952 1940
rect 12752 1792 12952 1802
rect 13432 1618 13931 1684
rect 10106 1210 11386 1410
rect 11244 356 11388 820
rect 12768 764 12832 1152
rect 12768 702 12832 712
rect 11776 552 11908 562
rect 11776 476 11908 486
rect 11244 346 11390 356
rect 11244 202 11246 346
rect 11244 192 11390 202
rect 9254 138 9322 186
rect 12352 171 12498 668
rect 12346 138 12498 171
rect 9254 59 12498 138
rect 13434 137 13500 1278
rect 13865 139 13931 1618
rect 14052 1416 14252 2306
rect 15360 1906 15520 1916
rect 15360 1812 15520 1822
rect 16888 1906 17048 1916
rect 16888 1812 17048 1822
rect 17548 1618 17740 1684
rect 14052 1216 15506 1416
rect 14030 996 14110 1006
rect 14110 916 16582 996
rect 14030 906 14110 916
rect 15364 346 15508 819
rect 16502 589 16582 916
rect 16888 762 16956 1108
rect 16952 730 16956 762
rect 16888 700 16952 710
rect 15890 554 16026 564
rect 15890 472 16026 482
rect 15506 200 15508 346
rect 15364 190 15506 200
rect 13353 -263 13753 137
rect 13831 130 14231 139
rect 17552 130 17616 1280
rect 13831 66 17616 130
rect 13831 -261 14231 66
rect 13677 -291 13743 -263
rect 17674 -291 17740 1618
rect 13677 -357 17740 -291
rect 2500 -834 2900 -672
rect 2500 -904 2526 -834
rect 2856 -904 2900 -834
rect 2500 -1072 2900 -904
<< via2 >>
rect 350 1612 606 1868
rect 7478 1704 7572 1804
rect 11218 1802 11418 1930
rect 12752 1802 12952 1930
rect 11776 486 11908 552
rect 15360 1822 15520 1906
rect 16888 1822 17048 1906
rect 15890 482 16026 554
<< metal3 >>
rect 11114 1930 17084 2016
rect 340 1868 616 1873
rect 340 1612 350 1868
rect 606 1866 616 1868
rect 11114 1866 11218 1930
rect 606 1804 11218 1866
rect 606 1704 7478 1804
rect 7572 1802 11218 1804
rect 11418 1802 12752 1930
rect 12952 1906 17084 1930
rect 12952 1822 15360 1906
rect 15520 1822 16888 1906
rect 17048 1822 17084 1906
rect 12952 1802 17084 1822
rect 7572 1760 17084 1802
rect 7572 1704 11370 1760
rect 606 1612 11370 1704
rect 340 1610 11370 1612
rect 340 1607 616 1610
rect 11764 557 11916 1760
rect 15880 559 16032 1760
rect 11764 552 11918 557
rect 11764 486 11776 552
rect 11908 486 11918 552
rect 11764 482 11918 486
rect 11766 481 11918 482
rect 15880 554 16036 559
rect 15880 482 15890 554
rect 16026 482 16036 554
rect 15880 477 16036 482
rect 15880 474 16032 477
use sky130_fd_bs_flash__special_sonosfet_star_EA7MKQ  X1
timestamp 1739996772
transform 1 0 4518 0 1 2482
box -519 -553 519 553
use charge_pump_neg_nmos  x2 ../charge_pump_neg_nmos
timestamp 1739484054
transform 1 0 5137 0 1 5264
box -4288 -1488 12990 4458
use charge_pump  x3 ../charge_pump
timestamp 1739252499
transform 1 0 5136 0 1 11293
box -4288 -1488 12990 4458
use vprog_controller  x4 ../vprog_controller
timestamp 1740594681
transform 1 0 9076 0 -1 -914
box 1324 -4282 4846 -1260
use inverter  x5 ../inverter
timestamp 1739087840
transform 1 0 7955 0 1 2357
box 0 -620 992 638
use inverter  x6
timestamp 1739087840
transform 1 0 851 0 1 1177
box 0 -620 992 638
use vprog_controller  x7
timestamp 1740594681
transform 1 0 13196 0 -1 -915
box 1324 -4282 4846 -1260
use sky130_fd_pr__pfet_g5v0d10v5_VPAE37  XM1
timestamp 1739996415
transform 1 0 10090 0 1 -873
box -2258 -347 2258 347
use sky130_fd_pr__pfet_g5v0d10v5_VPAE37  XM2
timestamp 1739996415
transform 1 0 5174 0 1 -873
box -2258 -347 2258 347
use sky130_fd_pr__pfet_g5v0d10v5_GJ3XY6  XM3
timestamp 1739996415
transform 1 0 1258 0 1 -873
box -1258 -347 1258 347
use sky130_fd_pr__pfet_g5v0d10v5_VPAE37  XM4
timestamp 1739996415
transform 1 0 6568 0 1 221
box -2258 -347 2258 347
use sky130_fd_pr__nfet_g5v0d10v5_9UU773  XM5
timestamp 1739996415
transform 1 0 6558 0 1 2484
box -278 -758 278 758
use sky130_fd_pr__nfet_g5v0d10v5_HQS8YU  XM8
timestamp 1739996415
transform 1 0 2601 0 1 2531
box -278 -458 278 458
<< labels >>
flabel metal2 -37 1529 363 1929 1 FreeSans 400 0 0 0 VDPWR
port 29 nsew signal output
flabel metal2 -103 9640 297 10040 1 FreeSans 400 0 0 0 VAPWR
port 30 nsew signal output
flabel metal2 -12 3096 388 3496 1 FreeSans 400 0 0 0 VGND
port 31 nsew signal output
flabel metal2 -75 7364 325 7764 1 FreeSans 400 0 0 0 clk
port 32 nsew signal output
flabel metal2 13353 -263 13753 137 1 FreeSans 400 0 0 0 prog_en
port 34 nsew signal output
flabel metal2 13831 -261 14231 139 1 FreeSans 400 0 0 0 erase_en
port 35 nsew signal output
flabel metal2 8974 2184 9374 2584 1 FreeSans 400 0 0 0 data_out
port 37 nsew signal output
flabel metal2 -22 933 378 1333 1 FreeSans 400 0 0 0 read_en
port 36 nsew signal output
flabel metal2 2500 -1072 2900 -672 1 FreeSans 400 0 0 0 VPROGMON
port 38 nsew signal output
<< end >>
