magic
tech sky130A
magscale 1 2
timestamp 1738900598
<< dnwell >>
rect 1413 -4193 3461 -2899
<< nwell >>
rect 1436 -1868 3334 -1260
rect 3734 -1868 4486 -1426
rect 1436 -2810 4584 -2656
rect 1324 -2932 4584 -2810
rect 1324 -3106 4612 -2932
rect 1324 -3986 1620 -3106
rect 3254 -3528 4612 -3106
rect 3254 -3986 3550 -3528
rect 1324 -4282 3550 -3986
<< mvnmos >>
rect 1556 -2102 2156 -2002
rect 2324 -2102 2924 -2002
rect 3092 -2102 3692 -2002
rect 3860 -2102 4460 -2002
rect 1556 -2312 2156 -2212
rect 2324 -2312 2924 -2212
rect 3092 -2312 3692 -2212
rect 3860 -2312 4460 -2212
rect 1556 -2522 2156 -2422
rect 2324 -2522 2924 -2422
rect 3092 -2522 3692 -2422
rect 3860 -2522 4460 -2422
rect 2494 -3386 2694 -3286
rect 2862 -3386 3062 -3286
rect 1808 -3642 2408 -3542
rect 2466 -3642 3066 -3542
rect 1808 -3852 2408 -3752
rect 2466 -3852 3066 -3752
rect 3672 -3738 4272 -3638
rect 3672 -3948 4272 -3848
rect 3672 -4158 4272 -4058
<< mvpmos >>
rect 1556 -1592 2156 -1492
rect 2324 -1592 2424 -1492
rect 2482 -1592 2582 -1492
rect 2640 -1592 2740 -1492
rect 2798 -1592 2898 -1492
rect 2956 -1592 3056 -1492
rect 3114 -1592 3214 -1492
rect 1556 -1802 2156 -1702
rect 2324 -1802 2424 -1702
rect 2482 -1802 2582 -1702
rect 2640 -1802 2740 -1702
rect 2798 -1802 2898 -1702
rect 2956 -1802 3056 -1702
rect 3114 -1802 3214 -1702
rect 3858 -1592 3958 -1492
rect 4016 -1592 4116 -1492
rect 4174 -1592 4274 -1492
rect 3858 -1802 3958 -1702
rect 4016 -1802 4116 -1702
rect 4174 -1802 4274 -1702
rect 1556 -2822 2156 -2722
rect 2324 -2822 2924 -2722
rect 3092 -2822 3692 -2722
rect 3860 -2822 4460 -2722
rect 3602 -3098 3702 -2998
rect 3760 -3098 3860 -2998
rect 3918 -3098 4018 -2998
rect 4076 -3098 4176 -2998
rect 4234 -3098 4334 -2998
rect 4392 -3098 4492 -2998
rect 3602 -3462 3702 -3362
rect 3760 -3462 3860 -3362
rect 3918 -3462 4018 -3362
rect 4076 -3462 4176 -3362
rect 4234 -3462 4334 -3362
rect 4392 -3462 4492 -3362
<< mvndiff >>
rect 1502 -2014 1556 -2002
rect 1502 -2090 1510 -2014
rect 1544 -2090 1556 -2014
rect 1502 -2102 1556 -2090
rect 2156 -2014 2324 -2002
rect 2156 -2090 2168 -2014
rect 2312 -2090 2324 -2014
rect 2156 -2102 2324 -2090
rect 2924 -2014 2978 -2002
rect 2924 -2090 2936 -2014
rect 2970 -2090 2978 -2014
rect 2924 -2102 2978 -2090
rect 3038 -2014 3092 -2002
rect 3038 -2090 3046 -2014
rect 3080 -2090 3092 -2014
rect 3038 -2102 3092 -2090
rect 3692 -2014 3860 -2002
rect 3692 -2090 3704 -2014
rect 3848 -2090 3860 -2014
rect 3692 -2102 3860 -2090
rect 4460 -2014 4514 -2002
rect 4460 -2090 4472 -2014
rect 4506 -2090 4514 -2014
rect 4460 -2102 4514 -2090
rect 1502 -2224 1556 -2212
rect 1502 -2300 1510 -2224
rect 1544 -2300 1556 -2224
rect 1502 -2312 1556 -2300
rect 2156 -2224 2324 -2212
rect 2156 -2300 2168 -2224
rect 2312 -2300 2324 -2224
rect 2156 -2312 2324 -2300
rect 2924 -2224 2978 -2212
rect 2924 -2300 2936 -2224
rect 2970 -2300 2978 -2224
rect 2924 -2312 2978 -2300
rect 3038 -2224 3092 -2212
rect 3038 -2300 3046 -2224
rect 3080 -2300 3092 -2224
rect 3038 -2312 3092 -2300
rect 3692 -2224 3860 -2212
rect 3692 -2300 3704 -2224
rect 3848 -2300 3860 -2224
rect 3692 -2312 3860 -2300
rect 4460 -2224 4514 -2212
rect 4460 -2300 4472 -2224
rect 4506 -2300 4514 -2224
rect 4460 -2312 4514 -2300
rect 1502 -2434 1556 -2422
rect 1502 -2510 1510 -2434
rect 1544 -2510 1556 -2434
rect 1502 -2522 1556 -2510
rect 2156 -2434 2324 -2422
rect 2156 -2510 2168 -2434
rect 2312 -2510 2324 -2434
rect 2156 -2522 2324 -2510
rect 2924 -2434 2978 -2422
rect 2924 -2510 2936 -2434
rect 2970 -2510 2978 -2434
rect 2924 -2522 2978 -2510
rect 3038 -2434 3092 -2422
rect 3038 -2510 3046 -2434
rect 3080 -2510 3092 -2434
rect 3038 -2522 3092 -2510
rect 3692 -2434 3860 -2422
rect 3692 -2510 3704 -2434
rect 3848 -2510 3860 -2434
rect 3692 -2522 3860 -2510
rect 4460 -2434 4514 -2422
rect 4460 -2510 4472 -2434
rect 4506 -2510 4514 -2434
rect 4460 -2522 4514 -2510
rect 2436 -3298 2494 -3286
rect 2436 -3374 2448 -3298
rect 2482 -3374 2494 -3298
rect 2436 -3386 2494 -3374
rect 2694 -3298 2862 -3286
rect 2694 -3374 2706 -3298
rect 2850 -3374 2862 -3298
rect 2694 -3386 2862 -3374
rect 3062 -3298 3120 -3286
rect 3062 -3374 3074 -3298
rect 3108 -3374 3120 -3298
rect 3062 -3386 3120 -3374
rect 1754 -3554 1808 -3542
rect 1754 -3630 1762 -3554
rect 1796 -3630 1808 -3554
rect 1754 -3642 1808 -3630
rect 2408 -3554 2466 -3542
rect 2408 -3630 2420 -3554
rect 2454 -3630 2466 -3554
rect 2408 -3642 2466 -3630
rect 3066 -3554 3120 -3542
rect 3066 -3630 3078 -3554
rect 3112 -3630 3120 -3554
rect 3066 -3642 3120 -3630
rect 1754 -3764 1808 -3752
rect 1754 -3840 1762 -3764
rect 1796 -3840 1808 -3764
rect 1754 -3852 1808 -3840
rect 2408 -3764 2466 -3752
rect 2408 -3840 2420 -3764
rect 2454 -3840 2466 -3764
rect 2408 -3852 2466 -3840
rect 3066 -3764 3120 -3752
rect 3066 -3840 3078 -3764
rect 3112 -3840 3120 -3764
rect 3066 -3852 3120 -3840
rect 3618 -3650 3672 -3638
rect 3618 -3726 3626 -3650
rect 3660 -3726 3672 -3650
rect 3618 -3738 3672 -3726
rect 4272 -3650 4326 -3638
rect 4272 -3726 4284 -3650
rect 4318 -3726 4326 -3650
rect 4272 -3738 4326 -3726
rect 3618 -3860 3672 -3848
rect 3618 -3936 3626 -3860
rect 3660 -3936 3672 -3860
rect 3618 -3948 3672 -3936
rect 4272 -3860 4326 -3848
rect 4272 -3936 4284 -3860
rect 4318 -3936 4326 -3860
rect 4272 -3948 4326 -3936
rect 3618 -4070 3672 -4058
rect 3618 -4146 3626 -4070
rect 3660 -4146 3672 -4070
rect 3618 -4158 3672 -4146
rect 4272 -4070 4326 -4058
rect 4272 -4146 4284 -4070
rect 4318 -4146 4326 -4070
rect 4272 -4158 4326 -4146
<< mvpdiff >>
rect 1502 -1504 1556 -1492
rect 1502 -1580 1510 -1504
rect 1544 -1580 1556 -1504
rect 1502 -1592 1556 -1580
rect 2156 -1504 2210 -1492
rect 2156 -1580 2168 -1504
rect 2202 -1580 2210 -1504
rect 2156 -1592 2210 -1580
rect 2270 -1504 2324 -1492
rect 2270 -1580 2278 -1504
rect 2312 -1580 2324 -1504
rect 2270 -1592 2324 -1580
rect 2424 -1504 2482 -1492
rect 2424 -1580 2436 -1504
rect 2470 -1580 2482 -1504
rect 2424 -1592 2482 -1580
rect 2582 -1504 2640 -1492
rect 2582 -1580 2594 -1504
rect 2628 -1580 2640 -1504
rect 2582 -1592 2640 -1580
rect 2740 -1504 2798 -1492
rect 2740 -1580 2752 -1504
rect 2786 -1580 2798 -1504
rect 2740 -1592 2798 -1580
rect 2898 -1504 2956 -1492
rect 2898 -1580 2910 -1504
rect 2944 -1580 2956 -1504
rect 2898 -1592 2956 -1580
rect 3056 -1504 3114 -1492
rect 3056 -1580 3068 -1504
rect 3102 -1580 3114 -1504
rect 3056 -1592 3114 -1580
rect 3214 -1504 3268 -1492
rect 3214 -1580 3226 -1504
rect 3260 -1580 3268 -1504
rect 3214 -1592 3268 -1580
rect 1502 -1714 1556 -1702
rect 1502 -1790 1510 -1714
rect 1544 -1790 1556 -1714
rect 1502 -1802 1556 -1790
rect 2156 -1714 2210 -1702
rect 2156 -1790 2168 -1714
rect 2202 -1790 2210 -1714
rect 2156 -1802 2210 -1790
rect 2270 -1714 2324 -1702
rect 2270 -1790 2278 -1714
rect 2312 -1790 2324 -1714
rect 2270 -1802 2324 -1790
rect 2424 -1714 2482 -1702
rect 2424 -1790 2436 -1714
rect 2470 -1790 2482 -1714
rect 2424 -1802 2482 -1790
rect 2582 -1714 2640 -1702
rect 2582 -1790 2594 -1714
rect 2628 -1790 2640 -1714
rect 2582 -1802 2640 -1790
rect 2740 -1714 2798 -1702
rect 2740 -1790 2752 -1714
rect 2786 -1790 2798 -1714
rect 2740 -1802 2798 -1790
rect 2898 -1714 2956 -1702
rect 2898 -1790 2910 -1714
rect 2944 -1790 2956 -1714
rect 2898 -1802 2956 -1790
rect 3056 -1714 3114 -1702
rect 3056 -1790 3068 -1714
rect 3102 -1790 3114 -1714
rect 3056 -1802 3114 -1790
rect 3214 -1714 3268 -1702
rect 3214 -1790 3226 -1714
rect 3260 -1790 3268 -1714
rect 3214 -1802 3268 -1790
rect 3800 -1504 3858 -1492
rect 3800 -1580 3812 -1504
rect 3846 -1580 3858 -1504
rect 3800 -1592 3858 -1580
rect 3958 -1504 4016 -1492
rect 3958 -1580 3970 -1504
rect 4004 -1580 4016 -1504
rect 3958 -1592 4016 -1580
rect 4116 -1504 4174 -1492
rect 4116 -1580 4128 -1504
rect 4162 -1580 4174 -1504
rect 4116 -1592 4174 -1580
rect 4274 -1504 4332 -1492
rect 4274 -1580 4286 -1504
rect 4320 -1580 4332 -1504
rect 4274 -1592 4332 -1580
rect 3800 -1714 3858 -1702
rect 3800 -1790 3812 -1714
rect 3846 -1790 3858 -1714
rect 3800 -1802 3858 -1790
rect 3958 -1714 4016 -1702
rect 3958 -1790 3970 -1714
rect 4004 -1790 4016 -1714
rect 3958 -1802 4016 -1790
rect 4116 -1714 4174 -1702
rect 4116 -1790 4128 -1714
rect 4162 -1790 4174 -1714
rect 4116 -1802 4174 -1790
rect 4274 -1714 4332 -1702
rect 4274 -1790 4286 -1714
rect 4320 -1790 4332 -1714
rect 4274 -1802 4332 -1790
rect 1502 -2734 1556 -2722
rect 1502 -2810 1510 -2734
rect 1544 -2810 1556 -2734
rect 1502 -2822 1556 -2810
rect 2156 -2734 2324 -2722
rect 2156 -2810 2168 -2734
rect 2312 -2810 2324 -2734
rect 2156 -2822 2324 -2810
rect 2924 -2734 2978 -2722
rect 2924 -2810 2936 -2734
rect 2970 -2810 2978 -2734
rect 2924 -2822 2978 -2810
rect 3038 -2734 3092 -2722
rect 3038 -2810 3046 -2734
rect 3080 -2810 3092 -2734
rect 3038 -2822 3092 -2810
rect 3692 -2734 3860 -2722
rect 3692 -2810 3704 -2734
rect 3848 -2810 3860 -2734
rect 3692 -2822 3860 -2810
rect 4460 -2734 4518 -2722
rect 4460 -2810 4472 -2734
rect 4506 -2810 4518 -2734
rect 4460 -2822 4518 -2810
rect 3548 -3010 3602 -2998
rect 3548 -3086 3556 -3010
rect 3590 -3086 3602 -3010
rect 3548 -3098 3602 -3086
rect 3702 -3010 3760 -2998
rect 3702 -3086 3714 -3010
rect 3748 -3086 3760 -3010
rect 3702 -3098 3760 -3086
rect 3860 -3010 3918 -2998
rect 3860 -3086 3872 -3010
rect 3906 -3086 3918 -3010
rect 3860 -3098 3918 -3086
rect 4018 -3010 4076 -2998
rect 4018 -3086 4030 -3010
rect 4064 -3086 4076 -3010
rect 4018 -3098 4076 -3086
rect 4176 -3010 4234 -2998
rect 4176 -3086 4188 -3010
rect 4222 -3086 4234 -3010
rect 4176 -3098 4234 -3086
rect 4334 -3010 4392 -2998
rect 4334 -3086 4346 -3010
rect 4380 -3086 4392 -3010
rect 4334 -3098 4392 -3086
rect 4492 -3010 4546 -2998
rect 4492 -3086 4504 -3010
rect 4538 -3086 4546 -3010
rect 4492 -3098 4546 -3086
rect 3548 -3374 3602 -3362
rect 3548 -3450 3556 -3374
rect 3590 -3450 3602 -3374
rect 3548 -3462 3602 -3450
rect 3702 -3374 3760 -3362
rect 3702 -3450 3714 -3374
rect 3748 -3450 3760 -3374
rect 3702 -3462 3760 -3450
rect 3860 -3374 3918 -3362
rect 3860 -3450 3872 -3374
rect 3906 -3450 3918 -3374
rect 3860 -3462 3918 -3450
rect 4018 -3374 4076 -3362
rect 4018 -3450 4030 -3374
rect 4064 -3450 4076 -3374
rect 4018 -3462 4076 -3450
rect 4176 -3374 4234 -3362
rect 4176 -3450 4188 -3374
rect 4222 -3450 4234 -3374
rect 4176 -3462 4234 -3450
rect 4334 -3374 4392 -3362
rect 4334 -3450 4346 -3374
rect 4380 -3450 4392 -3374
rect 4334 -3462 4392 -3450
rect 4492 -3374 4546 -3362
rect 4492 -3450 4504 -3374
rect 4538 -3450 4546 -3374
rect 4492 -3462 4546 -3450
<< mvndiffc >>
rect 1510 -2090 1544 -2014
rect 2168 -2090 2312 -2014
rect 2936 -2090 2970 -2014
rect 3046 -2090 3080 -2014
rect 3704 -2090 3848 -2014
rect 4472 -2090 4506 -2014
rect 1510 -2300 1544 -2224
rect 2168 -2300 2312 -2224
rect 2936 -2300 2970 -2224
rect 3046 -2300 3080 -2224
rect 3704 -2300 3848 -2224
rect 4472 -2300 4506 -2224
rect 1510 -2510 1544 -2434
rect 2168 -2510 2312 -2434
rect 2936 -2510 2970 -2434
rect 3046 -2510 3080 -2434
rect 3704 -2510 3848 -2434
rect 4472 -2510 4506 -2434
rect 2448 -3374 2482 -3298
rect 2706 -3374 2850 -3298
rect 3074 -3374 3108 -3298
rect 1762 -3630 1796 -3554
rect 2420 -3630 2454 -3554
rect 3078 -3630 3112 -3554
rect 1762 -3840 1796 -3764
rect 2420 -3840 2454 -3764
rect 3078 -3840 3112 -3764
rect 3626 -3726 3660 -3650
rect 4284 -3726 4318 -3650
rect 3626 -3936 3660 -3860
rect 4284 -3936 4318 -3860
rect 3626 -4146 3660 -4070
rect 4284 -4146 4318 -4070
<< mvpdiffc >>
rect 1510 -1580 1544 -1504
rect 2168 -1580 2202 -1504
rect 2278 -1580 2312 -1504
rect 2436 -1580 2470 -1504
rect 2594 -1580 2628 -1504
rect 2752 -1580 2786 -1504
rect 2910 -1580 2944 -1504
rect 3068 -1580 3102 -1504
rect 3226 -1580 3260 -1504
rect 1510 -1790 1544 -1714
rect 2168 -1790 2202 -1714
rect 2278 -1790 2312 -1714
rect 2436 -1790 2470 -1714
rect 2594 -1790 2628 -1714
rect 2752 -1790 2786 -1714
rect 2910 -1790 2944 -1714
rect 3068 -1790 3102 -1714
rect 3226 -1790 3260 -1714
rect 3812 -1580 3846 -1504
rect 3970 -1580 4004 -1504
rect 4128 -1580 4162 -1504
rect 4286 -1580 4320 -1504
rect 3812 -1790 3846 -1714
rect 3970 -1790 4004 -1714
rect 4128 -1790 4162 -1714
rect 4286 -1790 4320 -1714
rect 1510 -2810 1544 -2734
rect 2168 -2810 2312 -2734
rect 2936 -2810 2970 -2734
rect 3046 -2810 3080 -2734
rect 3704 -2810 3848 -2734
rect 4472 -2810 4506 -2734
rect 3556 -3086 3590 -3010
rect 3714 -3086 3748 -3010
rect 3872 -3086 3906 -3010
rect 4030 -3086 4064 -3010
rect 4188 -3086 4222 -3010
rect 4346 -3086 4380 -3010
rect 4504 -3086 4538 -3010
rect 3556 -3450 3590 -3374
rect 3714 -3450 3748 -3374
rect 3872 -3450 3906 -3374
rect 4030 -3450 4064 -3374
rect 4188 -3450 4222 -3374
rect 4346 -3450 4380 -3374
rect 4504 -3450 4538 -3374
<< mvpsubdiff >>
rect 3496 -1350 3530 -1326
rect 4612 -1350 4646 -1326
rect 3496 -1896 3530 -1872
rect 4612 -1908 4646 -1884
rect 1390 -1960 1424 -1936
rect 1390 -2588 1424 -2564
rect 1646 -3166 1706 -3132
rect 3168 -3166 3228 -3132
rect 1646 -3192 1680 -3166
rect 3194 -3192 3228 -3166
rect 1646 -3926 1680 -3900
rect 3194 -3926 3228 -3900
rect 1646 -3960 1706 -3926
rect 3168 -3960 3228 -3926
rect 4470 -3852 4768 -3828
rect 4470 -4102 4494 -3852
rect 4744 -4102 4768 -3852
rect 4470 -4126 4768 -4102
<< mvnsubdiff >>
rect 1530 -1360 1554 -1326
rect 3206 -1360 3230 -1326
rect 4386 -1516 4420 -1492
rect 4386 -1802 4420 -1778
rect 1390 -2910 1450 -2876
rect 3424 -2910 3484 -2876
rect 1390 -2936 1424 -2910
rect 3450 -2936 3484 -2910
rect 1390 -4182 1424 -4156
rect 3450 -4182 3484 -4156
rect 1390 -4216 1450 -4182
rect 3424 -4216 3484 -4182
<< mvpsubdiffcont >>
rect 3496 -1872 3530 -1350
rect 4612 -1884 4646 -1350
rect 1390 -2564 1424 -1960
rect 1706 -3166 3168 -3132
rect 1646 -3900 1680 -3192
rect 3194 -3900 3228 -3192
rect 1706 -3960 3168 -3926
rect 4494 -4102 4744 -3852
<< mvnsubdiffcont >>
rect 1554 -1360 3206 -1326
rect 4386 -1778 4420 -1516
rect 1450 -2910 3424 -2876
rect 1390 -4156 1424 -2936
rect 3450 -4156 3484 -2936
rect 1450 -4216 3424 -4182
<< poly >>
rect 1556 -1410 2156 -1394
rect 1556 -1444 1566 -1410
rect 2146 -1444 2156 -1410
rect 1556 -1492 2156 -1444
rect 2324 -1410 2424 -1394
rect 2324 -1444 2340 -1410
rect 2408 -1444 2424 -1410
rect 2324 -1492 2424 -1444
rect 2482 -1410 2582 -1394
rect 2482 -1444 2498 -1410
rect 2566 -1444 2582 -1410
rect 2482 -1492 2582 -1444
rect 2640 -1410 2740 -1394
rect 2640 -1444 2656 -1410
rect 2724 -1444 2740 -1410
rect 2640 -1492 2740 -1444
rect 2798 -1410 2898 -1394
rect 2798 -1444 2814 -1410
rect 2882 -1444 2898 -1410
rect 2798 -1492 2898 -1444
rect 2956 -1410 3056 -1394
rect 2956 -1444 2972 -1410
rect 3040 -1444 3056 -1410
rect 2956 -1492 3056 -1444
rect 3114 -1410 3214 -1394
rect 3114 -1444 3130 -1410
rect 3198 -1444 3214 -1410
rect 3114 -1492 3214 -1444
rect 1556 -1626 2156 -1592
rect 2324 -1626 2424 -1592
rect 2482 -1626 2582 -1592
rect 2640 -1626 2740 -1592
rect 2798 -1626 2898 -1592
rect 2956 -1626 3056 -1592
rect 3114 -1626 3214 -1592
rect 1556 -1702 2156 -1668
rect 2324 -1702 2424 -1668
rect 2482 -1702 2582 -1668
rect 2640 -1702 2740 -1668
rect 2798 -1702 2898 -1668
rect 2956 -1702 3056 -1668
rect 3114 -1702 3214 -1668
rect 1556 -1850 2156 -1802
rect 1556 -1884 1566 -1850
rect 2146 -1884 2156 -1850
rect 1556 -1900 2156 -1884
rect 2324 -1850 2424 -1802
rect 2324 -1884 2340 -1850
rect 2408 -1884 2424 -1850
rect 2324 -1900 2424 -1884
rect 2482 -1850 2582 -1802
rect 2482 -1884 2498 -1850
rect 2566 -1884 2582 -1850
rect 2482 -1900 2582 -1884
rect 2640 -1850 2740 -1802
rect 2640 -1884 2656 -1850
rect 2724 -1884 2740 -1850
rect 2640 -1900 2740 -1884
rect 2798 -1850 2898 -1802
rect 2798 -1884 2814 -1850
rect 2882 -1884 2898 -1850
rect 2798 -1900 2898 -1884
rect 2956 -1850 3056 -1802
rect 2956 -1884 2972 -1850
rect 3040 -1884 3056 -1850
rect 2956 -1900 3056 -1884
rect 3114 -1850 3214 -1802
rect 3114 -1884 3130 -1850
rect 3198 -1884 3214 -1850
rect 3114 -1900 3214 -1884
rect 3858 -1492 3958 -1464
rect 4016 -1492 4116 -1464
rect 4174 -1492 4274 -1464
rect 3858 -1702 3958 -1592
rect 4016 -1702 4116 -1592
rect 4174 -1702 4274 -1592
rect 3858 -1850 3958 -1802
rect 3858 -1884 3874 -1850
rect 3942 -1884 3958 -1850
rect 3858 -1900 3958 -1884
rect 4016 -1850 4116 -1802
rect 4016 -1884 4032 -1850
rect 4100 -1884 4116 -1850
rect 4016 -1900 4116 -1884
rect 4174 -1850 4274 -1802
rect 4174 -1884 4190 -1850
rect 4258 -1884 4274 -1850
rect 4174 -1900 4274 -1884
rect 1556 -2002 2156 -1968
rect 2324 -2002 2924 -1968
rect 3092 -2002 3692 -1968
rect 3860 -2002 4460 -1968
rect 1556 -2140 2156 -2102
rect 1556 -2174 1594 -2140
rect 2118 -2174 2156 -2140
rect 1556 -2212 2156 -2174
rect 2324 -2140 2924 -2102
rect 2324 -2174 2362 -2140
rect 2886 -2174 2924 -2140
rect 2324 -2212 2924 -2174
rect 3092 -2140 3692 -2102
rect 3092 -2174 3130 -2140
rect 3654 -2174 3692 -2140
rect 3092 -2212 3692 -2174
rect 3860 -2140 4460 -2102
rect 3860 -2174 3898 -2140
rect 4422 -2174 4460 -2140
rect 3860 -2212 4460 -2174
rect 1556 -2340 2156 -2312
rect 2324 -2340 2924 -2312
rect 3092 -2340 3692 -2312
rect 3860 -2340 4460 -2312
rect 1556 -2422 2156 -2390
rect 2324 -2422 2924 -2390
rect 3092 -2422 3692 -2390
rect 3860 -2422 4460 -2390
rect 1556 -2602 2156 -2522
rect 1556 -2642 1594 -2602
rect 2118 -2642 2156 -2602
rect 1556 -2722 2156 -2642
rect 2324 -2602 2924 -2522
rect 2324 -2642 2362 -2602
rect 2886 -2642 2924 -2602
rect 2324 -2722 2924 -2642
rect 3092 -2602 3692 -2522
rect 3092 -2642 3130 -2602
rect 3664 -2642 3692 -2602
rect 3092 -2722 3692 -2642
rect 3860 -2602 4460 -2522
rect 3860 -2642 3888 -2602
rect 4422 -2642 4460 -2602
rect 3860 -2722 4460 -2642
rect 1556 -2858 2156 -2822
rect 2324 -2858 2924 -2822
rect 3092 -2858 3692 -2822
rect 3860 -2858 4460 -2822
rect 2494 -3286 2694 -3198
rect 2862 -3214 3062 -3198
rect 2862 -3248 2878 -3214
rect 3046 -3248 3062 -3214
rect 2862 -3286 3062 -3248
rect 2494 -3424 2694 -3386
rect 2494 -3458 2510 -3424
rect 2678 -3458 2694 -3424
rect 2494 -3474 2694 -3458
rect 2862 -3474 3062 -3386
rect 1808 -3542 2408 -3516
rect 2466 -3542 3066 -3516
rect 1808 -3680 2408 -3642
rect 1808 -3714 1824 -3680
rect 2392 -3714 2408 -3680
rect 1808 -3752 2408 -3714
rect 2466 -3680 3066 -3642
rect 2466 -3714 2482 -3680
rect 3050 -3714 3066 -3680
rect 2466 -3752 3066 -3714
rect 1808 -3878 2408 -3852
rect 2466 -3878 3066 -3852
rect 3602 -2916 3702 -2900
rect 3602 -2950 3618 -2916
rect 3686 -2950 3702 -2916
rect 3602 -2998 3702 -2950
rect 3760 -2998 3860 -2900
rect 3918 -2998 4018 -2900
rect 4076 -2916 4176 -2900
rect 4076 -2950 4092 -2916
rect 4160 -2950 4176 -2916
rect 4076 -2998 4176 -2950
rect 4234 -2916 4334 -2900
rect 4234 -2950 4250 -2916
rect 4318 -2950 4334 -2916
rect 4234 -2998 4334 -2950
rect 4392 -2998 4492 -2900
rect 3602 -3196 3702 -3098
rect 3760 -3148 3860 -3098
rect 3760 -3182 3776 -3148
rect 3844 -3182 3860 -3148
rect 3760 -3196 3860 -3182
rect 3918 -3148 4018 -3098
rect 3918 -3182 3934 -3148
rect 4002 -3182 4018 -3148
rect 3918 -3196 4018 -3182
rect 4076 -3196 4176 -3098
rect 4234 -3196 4334 -3098
rect 4392 -3148 4492 -3098
rect 4392 -3182 4408 -3148
rect 4476 -3182 4492 -3148
rect 4392 -3196 4492 -3182
rect 3602 -3280 3702 -3264
rect 3602 -3314 3618 -3280
rect 3686 -3314 3702 -3280
rect 3602 -3362 3702 -3314
rect 3760 -3362 3860 -3264
rect 3918 -3362 4018 -3264
rect 4076 -3280 4176 -3264
rect 4076 -3314 4092 -3280
rect 4160 -3314 4176 -3280
rect 4076 -3362 4176 -3314
rect 4234 -3280 4334 -3264
rect 4234 -3314 4250 -3280
rect 4318 -3314 4334 -3280
rect 4234 -3362 4334 -3314
rect 4392 -3362 4492 -3264
rect 3602 -3560 3702 -3462
rect 3760 -3510 3860 -3462
rect 3760 -3544 3776 -3510
rect 3844 -3544 3860 -3510
rect 3760 -3560 3860 -3544
rect 3918 -3510 4018 -3462
rect 3918 -3544 3934 -3510
rect 4002 -3544 4018 -3510
rect 3918 -3560 4018 -3544
rect 4076 -3560 4176 -3462
rect 4234 -3560 4334 -3462
rect 4392 -3510 4492 -3462
rect 4392 -3544 4408 -3510
rect 4476 -3544 4492 -3510
rect 4392 -3560 4492 -3544
rect 3672 -3638 4272 -3604
rect 3672 -3776 4272 -3738
rect 3672 -3810 3682 -3776
rect 4262 -3810 4272 -3776
rect 3672 -3848 4272 -3810
rect 3672 -3986 4272 -3948
rect 3672 -4020 3682 -3986
rect 4262 -4020 4272 -3986
rect 3672 -4058 4272 -4020
rect 3672 -4190 4272 -4158
<< polycont >>
rect 1566 -1444 2146 -1410
rect 2340 -1444 2408 -1410
rect 2498 -1444 2566 -1410
rect 2656 -1444 2724 -1410
rect 2814 -1444 2882 -1410
rect 2972 -1444 3040 -1410
rect 3130 -1444 3198 -1410
rect 1566 -1884 2146 -1850
rect 2340 -1884 2408 -1850
rect 2498 -1884 2566 -1850
rect 2656 -1884 2724 -1850
rect 2814 -1884 2882 -1850
rect 2972 -1884 3040 -1850
rect 3130 -1884 3198 -1850
rect 3874 -1884 3942 -1850
rect 4032 -1884 4100 -1850
rect 4190 -1884 4258 -1850
rect 1594 -2174 2118 -2140
rect 2362 -2174 2886 -2140
rect 3130 -2174 3654 -2140
rect 3898 -2174 4422 -2140
rect 1594 -2642 2118 -2602
rect 2362 -2642 2886 -2602
rect 3130 -2642 3664 -2602
rect 3888 -2642 4422 -2602
rect 2878 -3248 3046 -3214
rect 2510 -3458 2678 -3424
rect 1824 -3714 2392 -3680
rect 2482 -3714 3050 -3680
rect 3618 -2950 3686 -2916
rect 4092 -2950 4160 -2916
rect 4250 -2950 4318 -2916
rect 3776 -3182 3844 -3148
rect 3934 -3182 4002 -3148
rect 4408 -3182 4476 -3148
rect 3618 -3314 3686 -3280
rect 4092 -3314 4160 -3280
rect 4250 -3314 4318 -3280
rect 3776 -3544 3844 -3510
rect 3934 -3544 4002 -3510
rect 4408 -3544 4476 -3510
rect 3682 -3810 4262 -3776
rect 3682 -4020 4262 -3986
<< locali >>
rect 1538 -1360 1554 -1326
rect 3206 -1360 3222 -1326
rect 3496 -1332 4646 -1326
rect 3530 -1338 4646 -1332
rect 1566 -1410 2146 -1394
rect 1566 -1460 2146 -1444
rect 2340 -1410 2408 -1394
rect 2340 -1460 2408 -1444
rect 2498 -1410 2566 -1394
rect 2498 -1460 2566 -1444
rect 2656 -1410 2724 -1394
rect 2656 -1460 2724 -1444
rect 2814 -1410 2882 -1394
rect 2814 -1460 2882 -1444
rect 2972 -1410 3040 -1394
rect 2972 -1460 3040 -1444
rect 3130 -1410 3198 -1394
rect 3130 -1460 3198 -1444
rect 1494 -1580 1510 -1504
rect 1544 -1580 1590 -1504
rect 1636 -1580 1654 -1504
rect 2152 -1580 2168 -1504
rect 2202 -1580 2218 -1504
rect 2262 -1580 2278 -1504
rect 2312 -1580 2328 -1504
rect 2420 -1580 2436 -1504
rect 2470 -1580 2486 -1504
rect 2578 -1580 2594 -1504
rect 2628 -1580 2644 -1504
rect 2736 -1580 2752 -1504
rect 2786 -1580 2802 -1504
rect 2894 -1580 2910 -1504
rect 2944 -1580 2960 -1504
rect 3052 -1580 3068 -1504
rect 3102 -1580 3118 -1504
rect 3210 -1580 3226 -1504
rect 3260 -1580 3276 -1504
rect 2420 -1614 2486 -1580
rect 2736 -1614 2802 -1580
rect 3052 -1614 3118 -1580
rect 2420 -1680 3118 -1614
rect 2420 -1714 2486 -1680
rect 2736 -1714 2802 -1680
rect 3052 -1714 3118 -1680
rect 3530 -1360 4612 -1338
rect 4270 -1504 4420 -1500
rect 3796 -1580 3812 -1504
rect 3846 -1580 3862 -1504
rect 3954 -1580 3970 -1504
rect 4004 -1580 4020 -1504
rect 4112 -1580 4128 -1504
rect 4162 -1580 4178 -1504
rect 4270 -1580 4286 -1504
rect 4320 -1516 4420 -1504
rect 4320 -1580 4386 -1516
rect 1494 -1790 1510 -1714
rect 1544 -1790 1560 -1714
rect 2152 -1790 2168 -1714
rect 2202 -1790 2218 -1714
rect 2262 -1790 2278 -1714
rect 2312 -1790 2328 -1714
rect 2420 -1790 2436 -1714
rect 2470 -1790 2486 -1714
rect 2578 -1790 2594 -1714
rect 2628 -1790 2644 -1714
rect 2736 -1790 2752 -1714
rect 2786 -1790 2802 -1714
rect 2894 -1790 2910 -1714
rect 2944 -1790 2960 -1714
rect 3052 -1790 3068 -1714
rect 3102 -1790 3118 -1714
rect 3210 -1790 3226 -1714
rect 3260 -1790 3276 -1714
rect 1566 -1850 2202 -1834
rect 2146 -1884 2202 -1850
rect 2324 -1884 2340 -1850
rect 2408 -1884 2424 -1850
rect 2482 -1884 2498 -1850
rect 2566 -1884 2582 -1850
rect 2640 -1884 2656 -1850
rect 2724 -1884 2740 -1850
rect 2798 -1884 2814 -1850
rect 2882 -1884 2898 -1850
rect 2956 -1884 2972 -1850
rect 3040 -1884 3056 -1850
rect 3114 -1884 3130 -1850
rect 3198 -1884 3214 -1850
rect 3954 -1624 4020 -1580
rect 4270 -1624 4386 -1580
rect 3954 -1670 4386 -1624
rect 3954 -1714 4020 -1670
rect 4270 -1714 4386 -1670
rect 3796 -1790 3812 -1714
rect 3846 -1790 3862 -1714
rect 3954 -1790 3970 -1714
rect 4004 -1790 4020 -1714
rect 4112 -1790 4128 -1714
rect 4162 -1790 4178 -1714
rect 4270 -1790 4286 -1714
rect 4320 -1778 4386 -1714
rect 4320 -1790 4420 -1778
rect 4270 -1794 4420 -1790
rect 1566 -1900 2202 -1884
rect 3496 -1888 3530 -1872
rect 3858 -1884 3874 -1850
rect 3942 -1884 3958 -1850
rect 4016 -1884 4032 -1850
rect 4100 -1884 4116 -1850
rect 4174 -1884 4190 -1850
rect 4258 -1884 4274 -1850
rect 4612 -1900 4646 -1884
rect 2146 -1924 2202 -1900
rect 2146 -1930 2350 -1924
rect 1390 -1960 1424 -1944
rect 2146 -1974 2270 -1930
rect 2146 -1980 2350 -1974
rect 3030 -2014 3096 -2008
rect 1494 -2090 1510 -2014
rect 1544 -2090 1560 -2014
rect 2152 -2090 2168 -2014
rect 2312 -2090 2328 -2014
rect 2920 -2090 2936 -2014
rect 2970 -2090 2986 -2014
rect 3030 -2090 3046 -2014
rect 3080 -2090 3096 -2014
rect 3688 -2090 3704 -2014
rect 3848 -2090 3864 -2014
rect 4456 -2090 4472 -2014
rect 4506 -2090 4522 -2014
rect 1594 -2140 2118 -2124
rect 1594 -2190 2118 -2174
rect 2362 -2140 2886 -2124
rect 2362 -2190 2886 -2174
rect 3130 -2140 3654 -2124
rect 3130 -2190 3654 -2174
rect 3898 -2140 4422 -2124
rect 3898 -2190 4422 -2174
rect 1494 -2300 1510 -2224
rect 1544 -2300 1560 -2224
rect 2152 -2300 2168 -2224
rect 2312 -2300 2328 -2224
rect 2920 -2300 2936 -2224
rect 2970 -2300 2986 -2224
rect 3030 -2300 3046 -2224
rect 3080 -2300 3096 -2224
rect 3688 -2300 3704 -2224
rect 3848 -2300 3864 -2224
rect 4456 -2300 4472 -2224
rect 4506 -2300 4522 -2224
rect 2710 -2340 3306 -2334
rect 2790 -2392 3226 -2340
rect 2710 -2398 3306 -2392
rect 1390 -2580 1424 -2564
rect 1494 -2510 1510 -2434
rect 1544 -2510 1560 -2434
rect 2152 -2510 2168 -2434
rect 2312 -2510 2328 -2434
rect 2920 -2510 2936 -2434
rect 2970 -2510 2986 -2434
rect 1494 -2586 1560 -2510
rect 1494 -2658 1504 -2586
rect 1550 -2658 1560 -2586
rect 1594 -2550 2118 -2544
rect 1594 -2596 1606 -2550
rect 2106 -2596 2118 -2550
rect 1594 -2602 2118 -2596
rect 1594 -2658 2118 -2642
rect 2362 -2550 2886 -2544
rect 2362 -2596 2374 -2550
rect 2874 -2596 2886 -2550
rect 2362 -2602 2886 -2596
rect 2362 -2658 2886 -2642
rect 2920 -2586 2986 -2510
rect 2920 -2658 2930 -2586
rect 2976 -2658 2986 -2586
rect 1494 -2734 1560 -2658
rect 2920 -2734 2986 -2658
rect 1494 -2810 1510 -2734
rect 1544 -2810 1560 -2734
rect 2152 -2810 2168 -2734
rect 2312 -2810 2328 -2734
rect 2920 -2810 2936 -2734
rect 2970 -2810 2986 -2734
rect 3030 -2510 3046 -2434
rect 3080 -2510 3096 -2434
rect 3688 -2510 3704 -2434
rect 3848 -2510 3864 -2434
rect 4456 -2510 4472 -2434
rect 4506 -2510 4522 -2434
rect 3030 -2586 3096 -2510
rect 3030 -2658 3040 -2586
rect 3086 -2658 3096 -2586
rect 3130 -2550 3664 -2544
rect 3130 -2596 3142 -2550
rect 3652 -2596 3664 -2550
rect 3130 -2602 3664 -2596
rect 3130 -2658 3664 -2642
rect 3888 -2550 4422 -2544
rect 3888 -2596 3900 -2550
rect 4410 -2596 4422 -2550
rect 3888 -2602 4422 -2596
rect 3888 -2658 4422 -2642
rect 4456 -2586 4522 -2510
rect 4456 -2658 4466 -2586
rect 4512 -2658 4522 -2586
rect 3030 -2734 3096 -2658
rect 4456 -2734 4522 -2658
rect 3030 -2810 3046 -2734
rect 3080 -2810 3096 -2734
rect 3688 -2810 3704 -2734
rect 3848 -2810 3864 -2734
rect 4456 -2810 4472 -2734
rect 4506 -2810 4522 -2734
rect 1390 -2910 1450 -2876
rect 3424 -2910 3484 -2876
rect 1390 -2936 1424 -2910
rect 3450 -2936 3484 -2910
rect 3286 -3012 3292 -2950
rect 3400 -3012 3406 -2950
rect 1646 -3166 1706 -3132
rect 3168 -3166 3228 -3132
rect 1646 -3192 1680 -3166
rect 2448 -3298 2482 -3282
rect 2690 -3298 2828 -3166
rect 3194 -3192 3228 -3166
rect 2862 -3248 2878 -3214
rect 3046 -3248 3062 -3214
rect 3074 -3298 3108 -3282
rect 2690 -3374 2706 -3298
rect 2850 -3374 2866 -3298
rect 2448 -3390 2482 -3374
rect 3074 -3390 3108 -3374
rect 2494 -3458 2510 -3424
rect 2678 -3458 2694 -3424
rect 1762 -3554 1796 -3538
rect 1762 -3646 1796 -3630
rect 2420 -3554 2454 -3538
rect 2420 -3646 2454 -3630
rect 3078 -3554 3112 -3538
rect 3078 -3646 3112 -3630
rect 1808 -3714 1824 -3680
rect 2392 -3714 2408 -3680
rect 2466 -3714 2482 -3680
rect 3050 -3714 3066 -3680
rect 1762 -3764 1796 -3748
rect 1762 -3856 1796 -3840
rect 2420 -3764 2454 -3748
rect 2420 -3856 2454 -3840
rect 3078 -3764 3112 -3748
rect 3078 -3856 3112 -3840
rect 1646 -3926 1680 -3900
rect 3286 -3454 3406 -3012
rect 3286 -3522 3292 -3454
rect 3400 -3522 3406 -3454
rect 3194 -3926 3228 -3900
rect 1646 -3960 1706 -3926
rect 3168 -3960 3228 -3926
rect 3556 -2916 4658 -2844
rect 3556 -2950 3618 -2916
rect 3686 -2950 4092 -2916
rect 4160 -2950 4250 -2916
rect 4318 -2950 4658 -2916
rect 3556 -2960 4658 -2950
rect 3556 -3010 3590 -2994
rect 3556 -3102 3590 -3086
rect 3714 -3010 3748 -2994
rect 3714 -3102 3748 -3086
rect 3872 -3010 3906 -2994
rect 3872 -3102 3906 -3086
rect 4030 -3010 4064 -2994
rect 4030 -3102 4064 -3086
rect 4188 -3010 4222 -2994
rect 4188 -3102 4222 -3086
rect 4346 -3010 4380 -2994
rect 4346 -3102 4380 -3086
rect 4504 -3010 4538 -2994
rect 4504 -3102 4538 -3086
rect 3602 -3182 3776 -3148
rect 3844 -3182 3934 -3148
rect 4002 -3182 4408 -3148
rect 4476 -3182 4492 -3148
rect 3602 -3212 4492 -3182
rect 3602 -3248 3614 -3212
rect 4480 -3248 4492 -3212
rect 3602 -3280 4492 -3248
rect 3602 -3314 3618 -3280
rect 3686 -3314 4092 -3280
rect 4160 -3314 4250 -3280
rect 4318 -3314 4492 -3280
rect 3556 -3374 3590 -3358
rect 3556 -3466 3590 -3450
rect 3714 -3374 3748 -3358
rect 3714 -3466 3748 -3450
rect 3872 -3374 3906 -3358
rect 3872 -3466 3906 -3450
rect 4030 -3374 4064 -3358
rect 4030 -3466 4064 -3450
rect 4188 -3374 4222 -3358
rect 4188 -3466 4222 -3450
rect 4346 -3374 4380 -3358
rect 4346 -3466 4380 -3450
rect 4504 -3374 4538 -3358
rect 4504 -3466 4538 -3450
rect 3556 -3510 4658 -3500
rect 3556 -3544 3776 -3510
rect 3844 -3544 3934 -3510
rect 4002 -3544 4408 -3510
rect 4476 -3544 4658 -3510
rect 3556 -3616 4658 -3544
rect 1390 -4182 1424 -4156
rect 3610 -3726 3626 -3650
rect 4268 -3726 4284 -3650
rect 4318 -3726 4334 -3650
rect 3682 -3776 4262 -3760
rect 3682 -3826 4262 -3810
rect 4478 -3852 4760 -3836
rect 3610 -3936 3626 -3860
rect 4268 -3936 4284 -3860
rect 4318 -3936 4334 -3860
rect 3682 -3986 4262 -3970
rect 3682 -4036 4262 -4020
rect 3610 -4146 3626 -4070
rect 4268 -4146 4284 -4070
rect 4318 -4146 4334 -4070
rect 4478 -4102 4494 -3852
rect 4744 -4102 4760 -3852
rect 4478 -4118 4760 -4102
rect 3450 -4182 3484 -4156
rect 1390 -4216 1450 -4182
rect 3424 -4216 3484 -4182
<< viali >>
rect 1554 -1360 3206 -1326
rect 3496 -1350 3530 -1332
rect 1572 -1444 2122 -1410
rect 2340 -1444 2408 -1410
rect 2498 -1444 2566 -1410
rect 2656 -1444 2724 -1410
rect 2814 -1444 2882 -1410
rect 2972 -1444 3040 -1410
rect 3130 -1444 3198 -1410
rect 1590 -1580 1636 -1504
rect 2168 -1580 2202 -1504
rect 2278 -1580 2312 -1504
rect 2594 -1580 2628 -1504
rect 2910 -1580 2944 -1504
rect 3226 -1580 3260 -1504
rect 3496 -1668 3530 -1350
rect 4612 -1350 4646 -1338
rect 3812 -1580 3846 -1504
rect 3970 -1580 4004 -1504
rect 4128 -1580 4162 -1504
rect 4286 -1580 4320 -1504
rect 1510 -1790 1544 -1714
rect 2168 -1790 2202 -1714
rect 2278 -1790 2312 -1714
rect 2594 -1790 2628 -1714
rect 2910 -1790 2944 -1714
rect 3226 -1790 3260 -1714
rect 1590 -1884 2140 -1850
rect 2340 -1884 2408 -1850
rect 2498 -1884 2566 -1850
rect 2656 -1884 2724 -1850
rect 2814 -1884 2882 -1850
rect 2972 -1884 3040 -1850
rect 3130 -1884 3198 -1850
rect 3812 -1790 3846 -1714
rect 3970 -1790 4004 -1714
rect 4128 -1790 4162 -1714
rect 4286 -1790 4320 -1714
rect 4386 -1778 4420 -1516
rect 4612 -1716 4646 -1350
rect 3874 -1884 3942 -1850
rect 4032 -1884 4100 -1850
rect 4190 -1884 4258 -1850
rect 1390 -2564 1424 -1960
rect 2270 -1974 2350 -1930
rect 1510 -2090 1544 -2014
rect 2168 -2090 2312 -2014
rect 2936 -2090 2970 -2014
rect 3046 -2090 3080 -2014
rect 3704 -2090 3848 -2014
rect 4472 -2090 4506 -2014
rect 1600 -2174 2112 -2140
rect 2368 -2174 2880 -2140
rect 3136 -2174 3648 -2140
rect 3904 -2174 4416 -2140
rect 1510 -2300 1544 -2224
rect 2168 -2300 2312 -2224
rect 2936 -2300 2970 -2224
rect 3046 -2300 3080 -2224
rect 3704 -2300 3848 -2224
rect 4472 -2300 4506 -2224
rect 1424 -2440 1442 -2388
rect 2710 -2392 2790 -2340
rect 3226 -2392 3306 -2340
rect 2168 -2510 2312 -2434
rect 1504 -2658 1550 -2586
rect 1606 -2596 2106 -2550
rect 2374 -2596 2874 -2550
rect 2930 -2658 2976 -2586
rect 2168 -2810 2312 -2734
rect 3704 -2510 3848 -2434
rect 3040 -2658 3086 -2586
rect 3142 -2596 3652 -2550
rect 3900 -2596 4410 -2550
rect 4466 -2658 4512 -2586
rect 3704 -2810 3848 -2734
rect 1450 -2910 2884 -2876
rect 3022 -2910 3424 -2876
rect 1390 -4154 1424 -2938
rect 3292 -3012 3400 -2950
rect 1706 -3166 2306 -3132
rect 2448 -3166 3166 -3132
rect 1646 -3898 1680 -3194
rect 2448 -3374 2482 -3298
rect 2878 -3248 3046 -3214
rect 2706 -3374 2850 -3298
rect 3074 -3374 3108 -3298
rect 2510 -3458 2678 -3424
rect 1762 -3630 1796 -3554
rect 2420 -3630 2454 -3554
rect 3078 -3630 3112 -3554
rect 1824 -3714 2374 -3680
rect 2500 -3714 3032 -3680
rect 1762 -3840 1796 -3764
rect 2420 -3840 2454 -3764
rect 3078 -3840 3112 -3764
rect 3194 -3898 3228 -3448
rect 3292 -3522 3400 -3454
rect 1706 -3960 2702 -3926
rect 2830 -3960 3168 -3926
rect 4658 -2960 4692 -2844
rect 3556 -3086 3590 -3010
rect 3714 -3080 3748 -3016
rect 3872 -3086 3906 -3010
rect 4030 -3080 4064 -3016
rect 4188 -3086 4222 -3010
rect 4346 -3080 4380 -3016
rect 4504 -3086 4538 -3010
rect 3614 -3248 4480 -3212
rect 3556 -3450 3590 -3374
rect 3714 -3444 3748 -3380
rect 3872 -3450 3906 -3374
rect 4030 -3444 4064 -3380
rect 4188 -3450 4222 -3374
rect 4346 -3444 4380 -3380
rect 4504 -3450 4538 -3374
rect 4658 -3616 4692 -3500
rect 3450 -4154 3484 -3656
rect 3626 -3726 3660 -3650
rect 3660 -3726 3702 -3650
rect 4284 -3726 4318 -3650
rect 3688 -3810 4256 -3776
rect 3626 -3936 3660 -3860
rect 3660 -3936 3702 -3860
rect 4284 -3936 4318 -3860
rect 3688 -4020 4256 -3986
rect 3626 -4146 3660 -4070
rect 3660 -4146 3702 -4070
rect 4284 -4146 4318 -4070
rect 4494 -4102 4744 -3852
rect 1450 -4216 3424 -4182
<< metal1 >>
rect 1542 -1326 3218 -1320
rect 1542 -1360 1554 -1326
rect 3206 -1360 3218 -1326
rect 1542 -1366 3218 -1360
rect 3490 -1332 4652 -1320
rect 1498 -1410 2128 -1398
rect 1498 -1444 1572 -1410
rect 2122 -1444 2128 -1410
rect 1498 -1456 2128 -1444
rect 1498 -1714 1556 -1456
rect 1498 -1790 1510 -1714
rect 1544 -1790 1556 -1714
rect 1498 -1924 1556 -1790
rect 1584 -1504 1642 -1492
rect 1584 -1580 1590 -1504
rect 1636 -1580 1642 -1504
rect 1584 -1838 1642 -1580
rect 2156 -1504 2214 -1366
rect 2328 -1410 3210 -1404
rect 2328 -1444 2340 -1410
rect 2408 -1444 2498 -1410
rect 2566 -1444 2656 -1410
rect 2724 -1444 2814 -1410
rect 2882 -1444 2972 -1410
rect 3040 -1444 3130 -1410
rect 3198 -1444 3210 -1410
rect 2328 -1450 3210 -1444
rect 2156 -1580 2168 -1504
rect 2202 -1580 2214 -1504
rect 2156 -1708 2214 -1580
rect 2266 -1504 3426 -1498
rect 2266 -1580 2278 -1504
rect 2312 -1580 2594 -1504
rect 2628 -1580 2910 -1504
rect 2944 -1580 3226 -1504
rect 3260 -1580 3276 -1504
rect 3420 -1580 3426 -1504
rect 2266 -1586 3426 -1580
rect 3338 -1708 3426 -1586
rect 3490 -1668 3496 -1332
rect 3530 -1338 4652 -1332
rect 3530 -1366 4612 -1338
rect 3530 -1668 3536 -1366
rect 3490 -1680 3536 -1668
rect 3800 -1504 3858 -1498
rect 3800 -1580 3812 -1504
rect 3846 -1580 3858 -1504
rect 3800 -1614 3858 -1580
rect 3958 -1504 4016 -1498
rect 3958 -1580 3970 -1504
rect 4004 -1580 4016 -1504
rect 3958 -1586 4016 -1580
rect 4116 -1504 4174 -1498
rect 4116 -1580 4128 -1504
rect 4162 -1580 4174 -1504
rect 4116 -1614 4174 -1580
rect 3800 -1680 4174 -1614
rect 3800 -1708 3858 -1680
rect 2156 -1714 3272 -1708
rect 2156 -1790 2168 -1714
rect 2312 -1790 2594 -1714
rect 2628 -1790 2910 -1714
rect 2944 -1790 3226 -1714
rect 3260 -1790 3272 -1714
rect 2156 -1796 3272 -1790
rect 3338 -1714 3858 -1708
rect 3338 -1790 3812 -1714
rect 3846 -1790 3858 -1714
rect 3338 -1796 3858 -1790
rect 3958 -1714 4016 -1708
rect 3958 -1790 3970 -1714
rect 4004 -1790 4016 -1714
rect 3958 -1796 4016 -1790
rect 4116 -1714 4174 -1680
rect 4116 -1790 4128 -1714
rect 4162 -1790 4174 -1714
rect 4116 -1796 4174 -1790
rect 4280 -1504 4426 -1492
rect 4280 -1580 4286 -1504
rect 4320 -1516 4426 -1504
rect 4320 -1580 4386 -1516
rect 4280 -1714 4386 -1580
rect 4280 -1790 4286 -1714
rect 4320 -1778 4386 -1714
rect 4420 -1756 4426 -1516
rect 4606 -1716 4612 -1366
rect 4646 -1716 4652 -1338
rect 4606 -1728 4652 -1716
rect 4420 -1778 4846 -1756
rect 4320 -1790 4846 -1778
rect 4280 -1802 4846 -1790
rect 1584 -1850 2146 -1838
rect 1584 -1884 1590 -1850
rect 2140 -1884 2146 -1850
rect 1584 -1896 2146 -1884
rect 2174 -1850 3284 -1834
rect 2174 -1884 2340 -1850
rect 2408 -1884 2498 -1850
rect 2566 -1884 2656 -1850
rect 2724 -1884 2814 -1850
rect 2882 -1884 2972 -1850
rect 3040 -1884 3130 -1850
rect 3198 -1884 3284 -1850
rect 2174 -1890 3284 -1884
rect 3862 -1850 4772 -1844
rect 3862 -1884 3874 -1850
rect 3942 -1884 4032 -1850
rect 4100 -1884 4190 -1850
rect 4258 -1884 4772 -1850
rect 3862 -1890 4772 -1884
rect 2174 -1924 2230 -1890
rect 3228 -1924 3284 -1890
rect 1384 -1960 1430 -1948
rect 1384 -2564 1390 -1960
rect 1424 -2376 1430 -1960
rect 1498 -1980 2230 -1924
rect 2258 -1930 3092 -1924
rect 2258 -1974 2270 -1930
rect 2350 -1974 3092 -1930
rect 2258 -1980 3092 -1974
rect 3228 -1980 4518 -1924
rect 1498 -2014 1556 -1980
rect 1498 -2090 1510 -2014
rect 1544 -2090 1556 -2014
rect 1498 -2224 1556 -2090
rect 2156 -2014 2324 -2008
rect 2156 -2090 2168 -2014
rect 2312 -2090 2324 -2014
rect 2156 -2096 2324 -2090
rect 2924 -2014 3092 -1980
rect 2924 -2090 2936 -2014
rect 2970 -2090 3046 -2014
rect 3080 -2090 3092 -2014
rect 1594 -2140 2118 -2128
rect 1594 -2174 1600 -2140
rect 2112 -2174 2118 -2140
rect 1594 -2186 2118 -2174
rect 2362 -2140 2886 -2128
rect 2362 -2174 2368 -2140
rect 2880 -2174 2886 -2140
rect 2362 -2186 2886 -2174
rect 1498 -2300 1510 -2224
rect 1544 -2300 1556 -2224
rect 1498 -2306 1556 -2300
rect 1810 -2334 1910 -2186
rect 2156 -2224 2324 -2218
rect 2156 -2300 2168 -2224
rect 2312 -2300 2324 -2224
rect 2156 -2306 2324 -2300
rect 1810 -2340 2802 -2334
rect 1424 -2388 1448 -2376
rect 1442 -2440 1448 -2388
rect 1424 -2452 1448 -2440
rect 1810 -2392 2710 -2340
rect 2790 -2392 2802 -2340
rect 1810 -2398 2802 -2392
rect 1424 -2564 1430 -2452
rect 1810 -2544 1910 -2398
rect 2156 -2434 2324 -2428
rect 2156 -2510 2168 -2434
rect 2312 -2510 2324 -2434
rect 2156 -2516 2324 -2510
rect 2572 -2544 2672 -2398
rect 2830 -2454 2886 -2186
rect 2924 -2224 3092 -2090
rect 3692 -2014 3860 -2008
rect 3692 -2090 3704 -2014
rect 3848 -2090 3860 -2014
rect 3692 -2096 3860 -2090
rect 4460 -2014 4518 -1980
rect 4460 -2090 4472 -2014
rect 4506 -2090 4518 -2014
rect 2924 -2300 2936 -2224
rect 2970 -2300 3046 -2224
rect 3080 -2300 3092 -2224
rect 2924 -2312 3092 -2300
rect 3130 -2140 3654 -2128
rect 3130 -2174 3136 -2140
rect 3648 -2174 3654 -2140
rect 3130 -2186 3654 -2174
rect 3898 -2130 4422 -2128
rect 3898 -2140 4364 -2130
rect 3898 -2174 3904 -2140
rect 3898 -2182 4364 -2174
rect 4416 -2182 4422 -2130
rect 3898 -2186 4422 -2182
rect 3130 -2454 3186 -2186
rect 3692 -2224 3860 -2218
rect 3692 -2300 3704 -2224
rect 3848 -2300 3860 -2224
rect 3692 -2306 3860 -2300
rect 4112 -2334 4212 -2186
rect 4460 -2224 4518 -2090
rect 4460 -2300 4472 -2224
rect 4506 -2300 4518 -2224
rect 4460 -2308 4518 -2300
rect 3214 -2340 4212 -2334
rect 3214 -2392 3226 -2340
rect 3306 -2392 4212 -2340
rect 3214 -2398 4212 -2392
rect 2830 -2510 3186 -2454
rect 3692 -2434 3860 -2428
rect 3692 -2510 3704 -2434
rect 3848 -2510 3860 -2434
rect 1384 -2576 1430 -2564
rect 1594 -2550 2886 -2544
rect 1498 -2586 1556 -2574
rect 1498 -2658 1504 -2586
rect 1550 -2654 1556 -2586
rect 1594 -2596 1606 -2550
rect 2106 -2596 2374 -2550
rect 2874 -2596 2886 -2550
rect 1594 -2602 2886 -2596
rect 2924 -2586 2982 -2510
rect 3692 -2516 3860 -2510
rect 4376 -2532 4698 -2498
rect 4358 -2538 4698 -2532
rect 4358 -2544 4364 -2538
rect 3130 -2550 4364 -2544
rect 4416 -2544 4698 -2538
rect 2924 -2654 2930 -2586
rect 1550 -2658 2930 -2654
rect 2976 -2658 2982 -2586
rect 1498 -2700 2982 -2658
rect 3034 -2586 3092 -2574
rect 3034 -2658 3040 -2586
rect 3086 -2654 3092 -2586
rect 3130 -2596 3142 -2550
rect 3652 -2596 3900 -2550
rect 4416 -2590 4422 -2544
rect 4410 -2596 4422 -2590
rect 3130 -2602 4422 -2596
rect 4460 -2586 4518 -2574
rect 4460 -2654 4466 -2586
rect 3086 -2658 4466 -2654
rect 4512 -2654 4518 -2586
rect 4512 -2658 4624 -2654
rect 3034 -2700 4624 -2658
rect 2156 -2734 2324 -2728
rect 2156 -2810 2168 -2734
rect 2312 -2810 2324 -2734
rect 2156 -2870 2324 -2810
rect 1384 -2876 2896 -2870
rect 1384 -2910 1450 -2876
rect 2884 -2910 2896 -2876
rect 1384 -2916 2896 -2910
rect 1384 -2938 1430 -2916
rect 1384 -4154 1390 -2938
rect 1424 -4154 1430 -2938
rect 2924 -2946 2982 -2700
rect 3692 -2734 3860 -2728
rect 3692 -2810 3704 -2734
rect 3848 -2810 3860 -2734
rect 3692 -2816 3860 -2810
rect 3010 -2876 3436 -2870
rect 3010 -2910 3022 -2876
rect 3424 -2910 3436 -2876
rect 3010 -2916 3436 -2910
rect 3280 -2946 3412 -2944
rect 2924 -2950 3412 -2946
rect 2924 -3012 3292 -2950
rect 3400 -3012 3412 -2950
rect 2924 -3016 3412 -3012
rect 3280 -3018 3412 -3016
rect 3462 -2976 4550 -2930
rect 3462 -3046 3508 -2976
rect 2340 -3092 3508 -3046
rect 3544 -3010 3602 -3004
rect 3544 -3086 3556 -3010
rect 3590 -3086 3602 -3010
rect 1634 -3132 2312 -3120
rect 1634 -3166 1706 -3132
rect 2306 -3166 2312 -3132
rect 1634 -3178 2312 -3166
rect 1634 -3194 1692 -3178
rect 1634 -3642 1646 -3194
rect 1610 -3656 1646 -3642
rect 1680 -3542 1692 -3194
rect 2340 -3418 2386 -3092
rect 3544 -3120 3602 -3086
rect 3702 -3016 3760 -3004
rect 3702 -3080 3704 -3016
rect 3756 -3080 3760 -3016
rect 3702 -3092 3760 -3080
rect 3860 -3010 3918 -2976
rect 3860 -3086 3872 -3010
rect 3906 -3086 3918 -3010
rect 3860 -3092 3918 -3086
rect 4018 -3016 4076 -3004
rect 4018 -3080 4020 -3016
rect 4072 -3080 4076 -3016
rect 4018 -3092 4076 -3080
rect 4176 -3010 4234 -3004
rect 4176 -3086 4188 -3010
rect 4222 -3086 4234 -3010
rect 4176 -3120 4234 -3086
rect 4334 -3016 4392 -3004
rect 4334 -3080 4336 -3016
rect 4388 -3080 4392 -3016
rect 4334 -3092 4392 -3080
rect 4492 -3010 4550 -2976
rect 4492 -3086 4504 -3010
rect 4538 -3086 4550 -3010
rect 4492 -3092 4550 -3086
rect 2442 -3132 3172 -3120
rect 2442 -3166 2448 -3132
rect 3166 -3166 3172 -3132
rect 2442 -3178 3172 -3166
rect 3518 -3166 4550 -3120
rect 3518 -3208 3564 -3166
rect 4578 -3194 4624 -2700
rect 2442 -3214 3564 -3208
rect 2442 -3248 2878 -3214
rect 3046 -3248 3564 -3214
rect 2442 -3254 3564 -3248
rect 2442 -3298 2488 -3254
rect 2442 -3374 2448 -3298
rect 2482 -3374 2488 -3298
rect 2442 -3386 2488 -3374
rect 2694 -3298 2862 -3292
rect 2694 -3374 2706 -3298
rect 2850 -3374 2862 -3298
rect 2694 -3380 2862 -3374
rect 3068 -3298 3114 -3286
rect 3068 -3374 3074 -3298
rect 3108 -3368 3114 -3298
rect 3518 -3294 3564 -3254
rect 3592 -3212 4624 -3194
rect 3592 -3248 3614 -3212
rect 4480 -3248 4624 -3212
rect 3592 -3266 4624 -3248
rect 4652 -2844 4698 -2544
rect 4652 -2960 4658 -2844
rect 4692 -2960 4698 -2844
rect 3518 -3340 4550 -3294
rect 3108 -3374 3508 -3368
rect 3068 -3414 3508 -3374
rect 3068 -3418 3114 -3414
rect 2340 -3424 3114 -3418
rect 2340 -3458 2510 -3424
rect 2678 -3458 3114 -3424
rect 2340 -3464 3114 -3458
rect 3182 -3448 3240 -3442
rect 1680 -3554 1802 -3542
rect 1680 -3630 1762 -3554
rect 1796 -3630 1802 -3554
rect 1680 -3642 1802 -3630
rect 1680 -3656 1754 -3642
rect 2340 -3674 2386 -3464
rect 1812 -3680 2386 -3674
rect 1812 -3714 1824 -3680
rect 2374 -3714 2386 -3680
rect 1812 -3720 2386 -3714
rect 2414 -3554 2460 -3538
rect 2414 -3630 2420 -3554
rect 2454 -3630 2460 -3554
rect 1610 -3752 1646 -3732
rect 1634 -3898 1646 -3752
rect 1680 -3752 1754 -3732
rect 1680 -3764 1802 -3752
rect 1680 -3840 1762 -3764
rect 1796 -3840 1802 -3764
rect 1680 -3852 1802 -3840
rect 2414 -3764 2460 -3630
rect 3072 -3554 3118 -3542
rect 2488 -3680 3044 -3674
rect 2488 -3714 2500 -3680
rect 3032 -3714 3044 -3680
rect 2488 -3720 3044 -3714
rect 2414 -3840 2420 -3764
rect 2454 -3840 2460 -3764
rect 1680 -3898 1692 -3852
rect 2414 -3856 2460 -3840
rect 1634 -3914 1692 -3898
rect 1634 -3926 2708 -3914
rect 1634 -3960 1706 -3926
rect 2702 -3960 2708 -3926
rect 1634 -3972 2708 -3960
rect 1384 -4176 1430 -4154
rect 2736 -4176 2796 -3720
rect 3072 -3840 3078 -3554
rect 3112 -3620 3118 -3554
rect 3112 -3626 3154 -3620
rect 3112 -3776 3154 -3770
rect 3112 -3840 3118 -3776
rect 3072 -3852 3118 -3840
rect 3182 -3898 3194 -3448
rect 3228 -3898 3240 -3448
rect 3286 -3454 3406 -3442
rect 3286 -3522 3292 -3454
rect 3400 -3522 3406 -3454
rect 3286 -3558 3406 -3522
rect 3462 -3484 3508 -3414
rect 3544 -3374 3602 -3368
rect 3544 -3450 3556 -3374
rect 3590 -3450 3602 -3374
rect 3544 -3484 3602 -3450
rect 3702 -3380 3760 -3368
rect 3702 -3444 3704 -3380
rect 3756 -3444 3760 -3380
rect 3702 -3456 3760 -3444
rect 3860 -3374 3918 -3340
rect 3860 -3450 3872 -3374
rect 3906 -3450 3918 -3374
rect 3860 -3456 3918 -3450
rect 4018 -3380 4076 -3368
rect 4018 -3444 4020 -3380
rect 4072 -3444 4076 -3380
rect 4018 -3456 4076 -3444
rect 4176 -3374 4234 -3368
rect 4176 -3450 4188 -3374
rect 4222 -3450 4234 -3374
rect 4176 -3484 4234 -3450
rect 4334 -3380 4392 -3368
rect 4334 -3444 4336 -3380
rect 4388 -3444 4392 -3380
rect 4334 -3456 4392 -3444
rect 4492 -3374 4550 -3340
rect 4492 -3450 4504 -3374
rect 4538 -3450 4550 -3374
rect 4492 -3456 4550 -3450
rect 3462 -3530 4590 -3484
rect 3286 -3616 3586 -3558
rect 3182 -3914 3240 -3898
rect 2824 -3926 3240 -3914
rect 2824 -3960 2830 -3926
rect 3168 -3960 3240 -3926
rect 2824 -3972 3240 -3960
rect 3444 -3656 3490 -3644
rect 3444 -4154 3450 -3656
rect 3484 -4154 3490 -3656
rect 3528 -3764 3586 -3616
rect 3620 -3650 3708 -3644
rect 4272 -3650 4388 -3644
rect 3614 -3726 3626 -3650
rect 3702 -3726 3714 -3650
rect 4272 -3726 4284 -3650
rect 4318 -3726 4388 -3650
rect 4544 -3656 4590 -3530
rect 4652 -3500 4698 -2960
rect 4652 -3616 4658 -3500
rect 4692 -3616 4698 -3500
rect 4652 -3628 4698 -3616
rect 4726 -3656 4772 -1890
rect 4544 -3702 4772 -3656
rect 3620 -3732 3708 -3726
rect 4272 -3730 4388 -3726
rect 4800 -3730 4846 -1802
rect 4272 -3732 4846 -3730
rect 3528 -3776 4262 -3764
rect 3528 -3810 3688 -3776
rect 4256 -3810 4262 -3776
rect 3528 -3822 4262 -3810
rect 4330 -3776 4846 -3732
rect 3528 -3974 3586 -3822
rect 4330 -3854 4388 -3776
rect 3620 -3860 3708 -3854
rect 4272 -3860 4388 -3854
rect 3614 -3936 3626 -3860
rect 3702 -3936 3714 -3860
rect 4272 -3936 4284 -3860
rect 4318 -3936 4388 -3860
rect 3620 -3942 3708 -3936
rect 4272 -3942 4388 -3936
rect 3528 -3986 4262 -3974
rect 3528 -4020 3688 -3986
rect 4256 -4020 4262 -3986
rect 3528 -4032 4262 -4020
rect 4330 -4064 4388 -3942
rect 3620 -4070 3708 -4064
rect 4272 -4070 4388 -4064
rect 3444 -4176 3490 -4154
rect 1384 -4182 3490 -4176
rect 1384 -4216 1450 -4182
rect 3424 -4216 3490 -4182
rect 1384 -4222 3490 -4216
rect 3614 -4146 3626 -4070
rect 3702 -4146 3714 -4070
rect 3614 -4180 3714 -4146
rect 4272 -4146 4284 -4070
rect 4318 -4146 4388 -4070
rect 4272 -4152 4388 -4146
rect 4482 -3852 4756 -3840
rect 4482 -4102 4494 -3852
rect 4744 -4102 4756 -3852
rect 4482 -4114 4756 -4102
rect 4482 -4180 4540 -4114
rect 3614 -4238 4540 -4180
<< via1 >>
rect 3276 -1580 3420 -1504
rect 2168 -1790 2202 -1714
rect 2202 -1790 2278 -1714
rect 2278 -1790 2312 -1714
rect 2168 -2090 2312 -2014
rect 2168 -2300 2312 -2224
rect 1390 -2440 1442 -2388
rect 2168 -2510 2312 -2434
rect 3704 -2090 3848 -2014
rect 4364 -2140 4416 -2130
rect 4364 -2174 4416 -2140
rect 4364 -2182 4416 -2174
rect 3704 -2300 3848 -2224
rect 3704 -2510 3848 -2434
rect 4364 -2550 4416 -2538
rect 4364 -2590 4410 -2550
rect 4410 -2590 4416 -2550
rect 2168 -2810 2312 -2734
rect 3704 -2810 3848 -2734
rect 3704 -3080 3714 -3016
rect 3714 -3080 3748 -3016
rect 3748 -3080 3756 -3016
rect 4020 -3080 4030 -3016
rect 4030 -3080 4064 -3016
rect 4064 -3080 4072 -3016
rect 4336 -3080 4346 -3016
rect 4346 -3080 4380 -3016
rect 4380 -3080 4388 -3016
rect 1610 -3732 1646 -3656
rect 1646 -3732 1680 -3656
rect 1680 -3732 1754 -3656
rect 3078 -3630 3112 -3626
rect 3112 -3630 3154 -3626
rect 3078 -3764 3154 -3630
rect 3078 -3770 3112 -3764
rect 3112 -3770 3154 -3764
rect 3704 -3444 3714 -3380
rect 3714 -3444 3748 -3380
rect 3748 -3444 3756 -3380
rect 4020 -3444 4030 -3380
rect 4030 -3444 4064 -3380
rect 4064 -3444 4072 -3380
rect 4336 -3444 4346 -3380
rect 4346 -3444 4380 -3380
rect 4380 -3444 4388 -3380
rect 3626 -3726 3702 -3650
rect 3626 -3936 3702 -3860
rect 3626 -4146 3702 -4070
rect 4494 -4102 4744 -3852
<< metal2 >>
rect 3270 -1580 3276 -1504
rect 3420 -1580 4022 -1504
rect 2162 -1790 2168 -1714
rect 2312 -1790 2318 -1714
rect 2168 -2014 3848 -2008
rect 2312 -2090 3704 -2014
rect 2168 -2224 3848 -2090
rect 2312 -2300 3704 -2224
rect 2168 -2382 3848 -2300
rect 1384 -2388 3848 -2382
rect 1384 -2440 1390 -2388
rect 1442 -2434 3848 -2388
rect 1442 -2440 2168 -2434
rect 1384 -2446 2168 -2440
rect 2312 -2510 3704 -2434
rect 2168 -2516 3848 -2510
rect 3946 -2602 4022 -1580
rect 4358 -2130 4422 -2124
rect 4358 -2182 4364 -2130
rect 4416 -2182 4422 -2130
rect 4358 -2188 4422 -2182
rect 4358 -2538 4422 -2532
rect 4358 -2590 4364 -2538
rect 4416 -2590 4422 -2538
rect 4358 -2596 4422 -2590
rect 3078 -2678 4022 -2602
rect 2168 -2734 2312 -2728
rect 2168 -2816 2312 -2810
rect 3078 -3626 3154 -2678
rect 3704 -2734 3848 -2728
rect 3704 -3010 3848 -2810
rect 3704 -3016 4388 -3010
rect 3756 -3080 4020 -3016
rect 4072 -3080 4336 -3016
rect 3704 -3380 4388 -3080
rect 3756 -3444 4020 -3380
rect 4072 -3444 4336 -3380
rect 3704 -3450 4388 -3444
rect 1610 -3656 1754 -3650
rect 1610 -3740 1754 -3732
rect 3078 -3776 3154 -3770
rect 3620 -3650 4750 -3644
rect 3620 -3726 3626 -3650
rect 3702 -3726 4750 -3650
rect 3620 -3852 4750 -3726
rect 3620 -3860 4494 -3852
rect 3620 -3936 3626 -3860
rect 3702 -3936 4494 -3860
rect 3620 -4070 4494 -3936
rect 3620 -4146 3626 -4070
rect 3702 -4102 4494 -4070
rect 4744 -4102 4750 -3852
rect 3702 -4146 4750 -4102
rect 3620 -4152 4750 -4146
<< labels >>
flabel viali 2168 -2510 2312 -2434 0 FreeMono 160 0 0 0 VGND
port 4 nsew
flabel viali 2168 -2090 2312 -2014 0 FreeMono 160 0 0 0 VGND
flabel viali 2936 -2300 2970 -2224 7 FreeMono 160 0 0 0 pos_mid
flabel viali 2936 -2090 2970 -2014 7 FreeMono 160 0 0 0 pos_mid
flabel viali 2168 -2300 2312 -2224 0 FreeMono 160 0 0 0 VGND
flabel viali 2168 -2810 2312 -2734 0 FreeMono 160 0 0 0 VDPWR
port 3 nsew
flabel locali 1494 -2810 1560 -2434 0 FreeMono 160 90 0 0 pos_en_b
flabel locali 2920 -2810 2986 -2434 0 FreeMono 160 90 0 0 pos_en_b
flabel locali 3030 -2810 3096 -2434 0 FreeMono 160 90 0 0 neg_en_b
flabel polycont 1594 -2174 2118 -2140 0 FreeMono 160 0 0 0 pos_en
flabel locali 1594 -2642 2118 -2602 0 FreeMono 160 0 0 0 pos_en
flabel polycont 2362 -2174 2886 -2140 0 FreeMono 160 0 0 0 pos_en_b
flabel locali 2362 -2642 2886 -2602 0 FreeMono 160 0 0 0 pos_en
flabel viali 1510 -2300 1544 -2224 3 FreeMono 160 0 0 0 pos_mid_b
flabel viali 1510 -2090 1544 -2014 3 FreeMono 160 0 0 0 pos_mid_b
flabel polycont 1566 -1444 2146 -1410 0 FreeMono 160 0 0 0 pos_mid_b
flabel viali 3130 -1884 3198 -1850 0 FreeMono 64 0 0 0 pos_mid_b
flabel viali 2972 -1884 3040 -1850 0 FreeMono 64 0 0 0 pos_mid_b
flabel viali 2814 -1884 2882 -1850 0 FreeMono 64 0 0 0 pos_mid_b
flabel viali 2656 -1884 2724 -1850 0 FreeMono 64 0 0 0 pos_mid_b
flabel viali 2498 -1884 2566 -1850 0 FreeMono 64 0 0 0 pos_mid_b
flabel viali 2340 -1884 2408 -1850 0 FreeMono 64 0 0 0 pos_mid_b
flabel viali 3226 -1580 3260 -1504 0 FreeMono 80 90 0 0 VOUT
flabel viali 2910 -1580 2944 -1504 0 FreeMono 80 90 0 0 VOUT
flabel viali 2594 -1580 2628 -1504 0 FreeMono 80 90 0 0 VOUT
flabel viali 2278 -1580 2312 -1504 0 FreeMono 80 90 0 0 VOUT
flabel locali 3068 -1580 3102 -1504 0 FreeMono 80 90 0 0 vintp
flabel locali 3068 -1790 3102 -1714 0 FreeMono 80 90 0 0 vintp
flabel locali 2752 -1580 2786 -1504 0 FreeMono 80 90 0 0 vintp
flabel locali 2752 -1790 2786 -1714 0 FreeMono 80 90 0 0 vintp
flabel locali 2436 -1580 2470 -1504 0 FreeMono 80 90 0 0 vintp
flabel locali 2436 -1790 2470 -1714 0 FreeMono 80 90 0 0 vintp
flabel viali 2340 -1444 2408 -1410 0 FreeMono 64 180 0 0 VDPWR
flabel viali 2498 -1444 2566 -1410 0 FreeMono 64 180 0 0 VDPWR
flabel viali 2656 -1444 2724 -1410 0 FreeMono 64 180 0 0 VDPWR
flabel viali 2814 -1444 2882 -1410 0 FreeMono 64 180 0 0 VDPWR
flabel viali 2972 -1444 3040 -1410 0 FreeMono 64 180 0 0 VDPWR
flabel viali 3130 -1444 3198 -1410 0 FreeMono 64 180 0 0 VDPWR
flabel polycont 1566 -1884 2146 -1850 0 FreeMono 160 180 0 0 pos_mid
flabel viali 1510 -1790 1544 -1714 3 FreeMono 160 0 0 0 pos_mid_b
flabel metal2 2168 -1790 2312 -1714 0 FreeMono 160 0 0 0 VPRGPOS
port 5 nsew
flabel viali 3226 -1790 3260 -1714 0 FreeMono 80 90 0 0 VPRGPOS
flabel viali 2910 -1790 2944 -1714 0 FreeMono 80 90 0 0 VPRGPOS
flabel viali 2594 -1790 2628 -1714 0 FreeMono 80 90 0 0 VPRGPOS
flabel viali 3078 -3840 3112 -3764 0 FreeMono 160 90 0 0 VOUT
flabel viali 3078 -3630 3112 -3554 0 FreeMono 160 90 0 0 VOUT
flabel polycont 2482 -3714 3050 -3680 0 FreeMono 160 0 0 0 VDPWR
flabel viali 2448 -3374 2482 -3298 0 FreeMono 64 90 0 0 neg_mid
flabel viali 2878 -3248 3046 -3214 0 FreeMono 160 0 0 0 neg_mid
flabel viali 2510 -3458 2678 -3424 0 FreeMono 160 0 0 0 neg_mid_b
flabel viali 3074 -3374 3108 -3298 0 FreeMono 64 90 0 0 neg_mid_b
flabel viali 2706 -3374 2850 -3298 0 FreeMono 160 0 0 0 VPRGNEG
flabel locali 3130 -2642 3664 -2602 0 FreeMono 160 0 0 0 neg_en
flabel viali 1390 -2278 1424 -2244 0 FreeMono 48 0 0 0 VGND
flabel viali 3556 -3086 3590 -3010 0 FreeMono 64 90 0 0 neg_mid
flabel viali 3556 -3450 3590 -3374 0 FreeMono 64 90 0 0 neg_mid_b
flabel locali 3618 -3314 3686 -3280 0 FreeMono 64 0 0 0 neg_en_b
flabel locali 3618 -2950 3686 -2916 0 FreeMono 64 0 0 0 neg_en
flabel locali 4408 -3544 4476 -3510 0 FreeMono 64 0 0 0 neg_en
flabel locali 3934 -3544 4002 -3510 0 FreeMono 64 0 0 0 neg_en
flabel locali 3776 -3544 3844 -3510 0 FreeMono 64 0 0 0 neg_en
flabel locali 4250 -2950 4318 -2916 0 FreeMono 64 0 0 0 neg_en
flabel locali 4092 -2950 4160 -2916 0 FreeMono 64 0 0 0 neg_en
flabel locali 4408 -3182 4476 -3148 0 FreeMono 64 0 0 0 neg_en_b
flabel locali 3934 -3182 4002 -3148 0 FreeMono 64 0 0 0 neg_en_b
flabel locali 3776 -3182 3844 -3148 0 FreeMono 64 0 0 0 neg_en_b
flabel locali 4250 -3314 4318 -3280 0 FreeMono 64 0 0 0 neg_en_b
flabel locali 4092 -3314 4160 -3280 0 FreeMono 64 0 0 0 neg_en_b
flabel mvpdiffc 3714 -3450 3748 -3374 0 FreeMono 64 90 0 0 VDPWR
flabel mvpdiffc 4030 -3450 4064 -3374 0 FreeMono 64 90 0 0 VDPWR
flabel viali 3872 -3450 3906 -3374 0 FreeMono 64 90 0 0 neg_mid
flabel viali 4188 -3450 4222 -3374 0 FreeMono 64 90 0 0 neg_mid_b
flabel mvpdiffc 4346 -3450 4380 -3374 0 FreeMono 64 90 0 0 VDPWR
flabel viali 4504 -3450 4538 -3374 0 FreeMono 64 90 0 0 neg_mid
flabel viali 4504 -3086 4538 -3010 0 FreeMono 64 90 0 0 neg_mid_b
flabel mvpdiffc 4346 -3086 4380 -3010 0 FreeMono 64 90 0 0 VDPWR
flabel viali 3872 -3086 3906 -3010 0 FreeMono 64 90 0 0 neg_mid_b
flabel viali 4188 -3086 4222 -3010 0 FreeMono 64 90 0 0 neg_mid
flabel mvpdiffc 4030 -3086 4064 -3010 0 FreeMono 64 90 0 0 VDPWR
flabel mvpdiffc 3714 -3086 3748 -3010 0 FreeMono 64 90 0 0 VDPWR
flabel locali 3888 -2642 4422 -2602 0 FreeMono 160 0 0 0 neg_en
flabel locali 4456 -2810 4522 -2434 0 FreeMono 160 90 0 0 neg_en_b
flabel viali 3704 -2810 3848 -2734 0 FreeMono 160 0 0 0 VDPWR
port 3 nsew
flabel viali 3704 -2090 3848 -2014 0 FreeMono 160 0 0 0 VGND
flabel viali 3704 -2300 3848 -2224 0 FreeMono 160 0 0 0 VGND
flabel viali 3704 -2510 3848 -2434 0 FreeMono 160 0 0 0 VGND
flabel viali 3046 -2090 3080 -2014 3 FreeMono 160 0 0 0 pos_mid
flabel viali 3046 -2300 3080 -2224 3 FreeMono 160 0 0 0 pos_mid
flabel viali 4472 -2090 4506 -2014 0 FreeMono 160 0 0 0 pos_mid_b
flabel viali 4472 -2300 4506 -2224 0 FreeMono 160 0 0 0 pos_mid_b
flabel polycont 3130 -2174 3654 -2140 0 FreeMono 160 0 0 0 pos_en_b
flabel polycont 3898 -2174 4422 -2140 0 FreeMono 160 0 0 0 pos_en
flabel viali 3626 -3726 3660 -3650 0 FreeMono 160 90 0 0 VGND
flabel viali 3626 -3936 3660 -3860 0 FreeMono 160 90 0 0 VGND
flabel viali 3626 -4146 3660 -4070 0 FreeMono 160 90 0 0 VGND
flabel polycont 3682 -3810 4262 -3776 0 FreeMono 160 180 0 0 pos_en_b
flabel polycont 3682 -4020 4262 -3986 0 FreeMono 160 180 0 0 pos_en_b
flabel viali 4284 -3726 4318 -3650 0 FreeMono 80 90 0 0 dcgint
flabel viali 4284 -3936 4318 -3860 0 FreeMono 80 90 0 0 dcgint
flabel viali 4284 -4146 4318 -4070 0 FreeMono 80 90 0 0 dcgint
flabel via1 4494 -4102 4744 -3852 0 FreeMono 160 0 0 0 VGND
port 4 nsew
flabel metal2 3078 -3770 3154 -3626 0 FreeMono 160 0 0 0 VOUT
flabel viali 4190 -1884 4258 -1850 0 FreeMono 64 0 0 0 neg_mid_b
flabel viali 4032 -1884 4100 -1850 0 FreeMono 64 0 0 0 neg_mid_b
flabel viali 3874 -1884 3942 -1850 0 FreeMono 64 0 0 0 neg_mid_b
rlabel viali 3812 -1580 3846 -1504 0 VOUT
rlabel viali 4128 -1580 4162 -1504 0 VOUT
rlabel viali 3812 -1790 3846 -1714 0 VOUT
rlabel viali 4128 -1790 4162 -1714 0 VOUT
flabel viali 4612 -1664 4646 -1630 0 FreeMono 48 0 0 0 VGND
flabel viali 3496 -1652 3530 -1618 0 FreeMono 48 0 0 0 VGND
flabel metal2 3276 -1580 3420 -1504 0 FreeMono 160 0 0 0 VOUT
port 2 nsew
flabel metal2 4358 -2188 4422 -2124 0 FreeMono 64 0 0 0 pos_en
port 0 nsew
flabel metal2 4358 -2596 4422 -2532 0 FreeMono 64 0 0 0 neg_en
port 1 nsew
flabel viali 2264 -1360 2298 -1326 0 FreeMono 48 0 0 0 VPRGPOS
flabel polycont 1824 -3714 2392 -3680 0 FreeMono 160 0 0 0 neg_mid_b
flabel viali 1762 -3630 1796 -3554 0 FreeMono 80 90 0 0 VPRGNEG
flabel metal2 1610 -3732 1754 -3656 0 FreeMono 160 0 0 0 VPRGNEG
port 6 nsew
flabel viali 1762 -3840 1796 -3764 0 FreeMono 80 90 0 0 VPRGNEG
<< end >>
