** sch_path: /home/amedcalf/projects/tt10-sonos-flash-party/xschem/charge_pump_tb.sch
**.subckt charge_pump_tb
V1 VAPWR GND 3.3
V2 CLK GND PULSE(0 1.8 0 0 0 250n 500n)
R1 ua[0] analog_pad 500 m=1
C1 ua[0] 0 2.5p m=1
C2 analog_pad 0 2.5p m=1
x1 VAPWR ua[0] CLK GND charge_pump
R2 ua[0] GND 10meg m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/amedcalf/open-asic/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt
.include ../../spice/charge_pump/pex/charge_pump.spice
*.include ../../spice/charge_pump/sch/charge_pump.spice




.tran 10n 100u
.save all
.options savecurrents

.control
run
write pump_tb.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VAPWR
.end
