magic
tech sky130A
magscale 1 2
timestamp 1740434279
<< error_s >>
rect 4496 2437 4540 2527
<< nwell >>
rect 3799 2745 5237 3235
rect 3799 2219 4289 2745
rect 4747 2219 5237 2745
rect 3799 1729 5237 2219
<< mvnsubdiff >>
rect 3999 1993 4087 2017
rect 3999 1953 4023 1993
rect 4063 1953 4087 1993
rect 3999 1929 4087 1953
<< mvnsubdiffcont >>
rect 4023 1953 4063 1993
<< locali >>
rect 4007 1993 4079 2009
rect 4007 1953 4023 1993
rect 4063 1953 4079 1993
rect 4007 1937 4079 1953
<< viali >>
rect 2368 2540 2406 2858
rect 6746 1874 6786 3092
<< metal1 >>
rect 12144 13506 12154 13518
rect 11706 13364 12154 13506
rect 12412 13506 12422 13518
rect 14248 13506 14392 13510
rect 12412 13364 14392 13506
rect 11706 13362 14392 13364
rect 3450 12528 5382 12728
rect 3450 9990 3650 12528
rect 3748 12027 3848 12042
rect 3748 11927 5284 12027
rect 3438 9984 3662 9990
rect 3438 9784 3450 9984
rect 3650 9784 3662 9984
rect 3438 9778 3662 9784
rect 3748 7690 3848 11927
rect 3931 9771 3941 9981
rect 4151 9771 5390 9981
rect 112 7590 122 7690
rect 222 7590 3848 7690
rect 3748 5998 3848 7590
rect 5180 6492 5390 9771
rect 3748 5898 5286 5998
rect 2340 3168 2350 3260
rect 2442 3168 2452 3260
rect 2350 2858 2442 3168
rect 6740 3092 6792 3104
rect 6532 3026 6672 3058
rect 2350 2540 2368 2858
rect 2406 2600 2442 2858
rect 2406 2540 2534 2600
rect 2350 2508 2534 2540
rect 2581 2298 2609 2801
rect 4462 2568 4472 2622
rect 4538 2568 4548 2622
rect 2666 2466 4466 2502
rect 4558 2458 6478 2498
rect 4460 2344 4470 2400
rect 4544 2344 4554 2400
rect 6640 2392 6672 3026
rect 6740 2392 6746 3092
rect 6640 2334 6746 2392
rect 2562 2072 2626 2298
rect 14 2010 2626 2072
rect 14 2008 2622 2010
rect 14 1214 78 2008
rect 6640 1946 6672 2334
rect 6568 1914 6672 1946
rect 6740 1874 6746 2334
rect 6786 2392 6792 3092
rect 6786 2334 8244 2392
rect 6786 1874 6792 2334
rect 6740 1862 6792 1874
rect 6746 1834 6792 1862
rect 116 1670 126 1790
rect 246 1670 578 1790
rect 458 1550 578 1670
rect 458 1430 1041 1550
rect 14 1150 274 1214
rect 338 1150 1379 1214
rect 1690 1150 3904 1214
rect 7261 1191 7319 2334
rect 8574 2330 8992 2394
rect 9056 2330 9066 2394
rect 682 896 1032 900
rect 682 844 692 896
rect 744 844 1032 896
rect 682 836 1032 844
rect 3840 146 3904 1150
rect 4149 1133 7319 1191
rect 4149 727 4207 1133
rect 4149 669 4553 727
rect 5726 146 5790 860
rect 14248 346 14392 13362
rect 11236 202 11246 346
rect 11390 202 15364 346
rect 15354 200 15364 202
rect 15506 202 15520 346
rect 15506 200 15516 202
rect 3840 82 5790 146
<< via1 >>
rect 12154 13364 12412 13518
rect 3450 9784 3650 9984
rect 3941 9771 4151 9981
rect 122 7590 222 7690
rect 2350 3168 2442 3260
rect 4472 2568 4538 2622
rect 4470 2344 4544 2400
rect 126 1670 246 1790
rect 274 1150 338 1214
rect 8992 2330 9056 2394
rect 692 844 744 896
rect 11246 202 11390 346
rect 15364 200 15506 346
<< metal2 >>
rect 11520 13518 12412 13542
rect 11520 13366 12154 13518
rect 12154 13354 12412 13364
rect 4802 11341 5572 11541
rect -103 9991 4114 10040
rect -103 9984 4151 9991
rect -103 9784 3450 9984
rect 3650 9981 4151 9984
rect 3650 9784 3941 9981
rect -103 9771 3941 9784
rect -103 9761 4151 9771
rect -103 9640 4114 9761
rect -75 7690 325 7764
rect -75 7590 122 7690
rect 222 7590 325 7690
rect -75 7364 325 7590
rect 4802 5512 5002 11341
rect 11536 7342 11929 7528
rect 4802 5312 5650 5512
rect -12 3464 3608 3496
rect 4802 3464 5002 5312
rect 11743 3733 11929 7342
rect -12 3264 5002 3464
rect 10679 3547 14957 3733
rect -12 3260 3608 3264
rect -12 3168 2350 3260
rect 2442 3168 3608 3260
rect -12 3096 3608 3168
rect -37 1790 363 1929
rect -37 1670 126 1790
rect 246 1670 363 1790
rect -37 1529 363 1670
rect -22 1214 378 1333
rect -22 1150 274 1214
rect 338 1150 378 1214
rect -22 933 378 1150
rect 680 896 754 3096
rect 10679 2739 10865 3547
rect 14771 2733 14957 3547
rect 4464 2632 4536 2634
rect 4464 2622 4538 2632
rect 4464 2568 4472 2622
rect 4464 2558 4538 2568
rect 4464 2410 4536 2558
rect 4464 2400 4544 2410
rect 4464 2344 4470 2400
rect 4464 2334 4544 2344
rect 8974 2394 9374 2584
rect 4464 1524 4536 2334
rect 8974 2330 8992 2394
rect 9056 2330 9374 2394
rect 8974 2184 9374 2330
rect 13432 1618 13931 1684
rect 17548 1618 17740 1684
rect 4464 1452 9326 1524
rect 680 844 692 896
rect 744 844 754 896
rect 680 834 754 844
rect 9254 186 9326 1452
rect 11244 356 11388 820
rect 11244 346 11390 356
rect 11244 202 11246 346
rect 11244 192 11390 202
rect 9254 138 9322 186
rect 12352 171 12498 668
rect 12346 138 12498 171
rect 9254 59 12498 138
rect 13434 137 13500 1278
rect 13865 139 13931 1618
rect 15364 346 15508 819
rect 15506 200 15508 346
rect 15364 190 15506 200
rect 13353 -263 13753 137
rect 13831 130 14231 139
rect 17552 130 17616 1280
rect 13831 66 17616 130
rect 13831 -261 14231 66
rect 13677 -291 13743 -263
rect 17674 -291 17740 1618
rect 13677 -357 17740 -291
use sky130_fd_bs_flash__special_sonosfet_star_EA7MKQ  X1
timestamp 1739996772
transform 1 0 4518 0 1 2482
box -519 -553 519 553
use charge_pump_neg_nmos  x2 ../charge_pump_neg_nmos
timestamp 1740420321
transform 1 0 5137 0 1 5264
box -4288 -1488 12990 4458
use charge_pump  x3 ../charge_pump
timestamp 1740420321
transform 1 0 5136 0 1 11293
box -4288 -1488 12990 4458
use vprog_controller  x4 ../vprog_controller
timestamp 1738900598
transform 1 0 9076 0 -1 -914
box 1324 -4282 4846 -1260
use inverter  x5 ../inverter
timestamp 1739087840
transform 1 0 7735 0 1 2357
box 0 -620 992 638
use inverter  x6
timestamp 1739087840
transform 1 0 851 0 1 1177
box 0 -620 992 638
use vprog_controller  x7
timestamp 1738900598
transform 1 0 13196 0 -1 -915
box 1324 -4282 4846 -1260
use sky130_fd_pr__pfet_g5v0d10v5_VPAE37  XM1
timestamp 1739996415
transform 1 0 10090 0 1 -873
box -2258 -347 2258 347
use sky130_fd_pr__pfet_g5v0d10v5_VPAE37  XM2
timestamp 1739996415
transform 1 0 5174 0 1 -873
box -2258 -347 2258 347
use sky130_fd_pr__pfet_g5v0d10v5_GJ3XY6  XM3
timestamp 1739996415
transform 1 0 1258 0 1 -873
box -1258 -347 1258 347
use sky130_fd_pr__pfet_g5v0d10v5_VPAE37  XM4
timestamp 1739996415
transform 1 0 6566 0 1 707
box -2258 -347 2258 347
use sky130_fd_pr__nfet_g5v0d10v5_9UU773  XM5
timestamp 1739996415
transform 1 0 6558 0 1 2484
box -278 -758 278 758
use sky130_fd_pr__nfet_g5v0d10v5_HQS8YU  XM8
timestamp 1739996415
transform 1 0 2601 0 1 2531
box -278 -458 278 458
<< labels >>
flabel metal2 -37 1529 363 1929 1 FreeSans 400 0 0 0 VDPWR
port 29 nsew signal output
flabel metal2 -103 9640 297 10040 1 FreeSans 400 0 0 0 VAPWR
port 30 nsew signal output
flabel metal2 -12 3096 388 3496 1 FreeSans 400 0 0 0 VGND
port 31 nsew signal output
flabel metal2 -75 7364 325 7764 1 FreeSans 400 0 0 0 clk
port 32 nsew signal output
flabel metal2 13353 -263 13753 137 1 FreeSans 400 0 0 0 prog_en
port 34 nsew signal output
flabel metal2 13831 -261 14231 139 1 FreeSans 400 0 0 0 erase_en
port 35 nsew signal output
flabel metal2 8974 2184 9374 2584 1 FreeSans 400 0 0 0 data_out
port 37 nsew signal output
flabel metal2 -22 933 378 1333 1 FreeSans 400 0 0 0 read_en
port 36 nsew signal output
<< end >>
