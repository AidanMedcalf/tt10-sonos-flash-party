* NGSPICE file created from vprog_controller.ext - technology: sky130A

.subckt vprog_controller pos_en neg_en VOUT VDPWR VGND VPRGPOS VPRGNEG
X0 VDPWR neg_en neg_mid VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X1 pos_mid_b pos_en VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X2 VOUT neg_mid_b dcgint dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X3 VDPWR pos_en pos_en_b VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X4 VOUT VDPWR vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X5 dcgint neg_mid_b VOUT dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X6 pos_mid_b pos_en VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X7 vintp pos_mid_b VPRGPOS VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X8 neg_en_b neg_en VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X9 VPRGPOS pos_mid_b vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X10 VOUT neg_mid_b dcgint dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X11 dcgint neg_mid_b VOUT dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X12 pos_mid pos_en_b VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X13 neg_en_b neg_en VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=3
X14 neg_mid neg_en VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X15 vintp pos_mid_b VPRGPOS VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X16 VDPWR neg_en_b neg_mid_b VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X17 VDPWR neg_en_b neg_mid_b VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X18 a_2408_n3852# neg_mid_b VPRGNEG VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X19 VDPWR neg_en_b neg_mid_b VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X20 neg_mid neg_en VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X21 vintp VDPWR VOUT VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X22 pos_mid pos_en_b VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X23 neg_mid neg_en VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X24 VOUT VDPWR vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X25 VGND pos_en_b pos_mid VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X26 pos_en_b pos_en VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X27 a_2408_n3852# neg_mid_b VPRGNEG VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X28 vintp VDPWR VOUT VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X29 VGND pos_en_b pos_mid VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X30 pos_en_b pos_en VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X31 VPRGPOS pos_mid_b vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X32 VGND neg_en neg_en_b VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X33 vintp pos_mid_b VPRGPOS VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X34 dcgint pos_en_b VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X35 VDPWR neg_en neg_mid VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X36 VDPWR neg_en neg_en_b VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X37 VDPWR neg_en neg_mid VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X38 dcgint pos_en_b VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X39 VPRGPOS pos_mid pos_mid_b VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X40 neg_mid_b neg_mid VPRGNEG VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=1
X41 neg_mid_b neg_en_b VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X42 neg_mid_b neg_en_b VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X43 VOUT VDPWR vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X44 VPRGNEG neg_mid_b neg_mid VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.145 ps=1.58 w=0.5 l=1
X45 dcgint neg_mid_b VOUT dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X46 vintp VDPWR VOUT VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X47 VGND pos_en pos_mid_b VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X48 VOUT VDPWR a_2408_n3852# VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X49 dcgint pos_en_b VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X50 VPRGPOS pos_mid_b pos_mid VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X51 VGND pos_en pos_mid_b VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X52 VOUT VDPWR a_2408_n3852# VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X53 VPRGPOS pos_mid_b vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X54 neg_mid_b neg_en_b VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X55 dcgint neg_mid_b VOUT dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X56 VGND pos_en pos_en_b VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
.ends

