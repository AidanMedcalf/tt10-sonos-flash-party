magic
tech sky130A
magscale 1 2
timestamp 1739484054
<< dnwell >>
rect 877 1613 1831 2723
rect 3091 1613 4045 2723
rect 5305 1613 6259 2723
<< nwell >>
rect 768 2516 1940 2832
rect 768 1820 1084 2516
rect 1624 1820 1940 2516
rect 768 1504 1940 1820
rect 2982 2516 4154 2832
rect 2982 1820 3298 2516
rect 3838 1820 4154 2516
rect 2982 1504 4154 1820
rect 5196 2516 6368 2832
rect 5196 1820 5512 2516
rect 6052 1820 6368 2516
rect 5196 1504 6368 1820
rect -24 694 1940 1504
<< pwell >>
rect 1084 1820 1624 2516
rect 3298 1820 3838 2516
rect 5512 1820 6052 2516
rect 6 12 1910 608
<< mvnmos >>
rect 1304 2068 1404 2268
rect 3518 2068 3618 2268
rect 5732 2068 5832 2268
rect 234 370 434 470
rect 650 370 850 470
rect 1066 270 1266 470
rect 1482 270 1682 470
<< mvpmos >>
rect 234 906 434 1006
rect 650 906 850 1006
rect 1066 906 1266 1206
rect 1482 906 1682 1206
<< mvndiff >>
rect 1246 2256 1304 2268
rect 1246 2080 1258 2256
rect 1292 2080 1304 2256
rect 1246 2068 1304 2080
rect 1404 2256 1462 2268
rect 1404 2080 1416 2256
rect 1450 2080 1462 2256
rect 1404 2068 1462 2080
rect 3460 2256 3518 2268
rect 3460 2080 3472 2256
rect 3506 2080 3518 2256
rect 3460 2068 3518 2080
rect 3618 2256 3676 2268
rect 3618 2080 3630 2256
rect 3664 2080 3676 2256
rect 3618 2068 3676 2080
rect 5674 2256 5732 2268
rect 5674 2080 5686 2256
rect 5720 2080 5732 2256
rect 5674 2068 5732 2080
rect 5832 2256 5890 2268
rect 5832 2080 5844 2256
rect 5878 2080 5890 2256
rect 5832 2068 5890 2080
rect 176 458 234 470
rect 176 382 188 458
rect 222 382 234 458
rect 176 370 234 382
rect 434 458 492 470
rect 434 382 446 458
rect 480 382 492 458
rect 434 370 492 382
rect 592 458 650 470
rect 592 382 604 458
rect 638 382 650 458
rect 592 370 650 382
rect 850 458 908 470
rect 850 382 862 458
rect 896 382 908 458
rect 850 370 908 382
rect 1008 458 1066 470
rect 1008 282 1020 458
rect 1054 282 1066 458
rect 1008 270 1066 282
rect 1266 458 1324 470
rect 1266 282 1278 458
rect 1312 282 1324 458
rect 1266 270 1324 282
rect 1424 458 1482 470
rect 1424 282 1436 458
rect 1470 282 1482 458
rect 1424 270 1482 282
rect 1682 458 1740 470
rect 1682 282 1694 458
rect 1728 282 1740 458
rect 1682 270 1740 282
<< mvpdiff >>
rect 1008 1194 1066 1206
rect 176 994 234 1006
rect 176 918 188 994
rect 222 918 234 994
rect 176 906 234 918
rect 434 994 492 1006
rect 434 918 446 994
rect 480 918 492 994
rect 434 906 492 918
rect 592 994 650 1006
rect 592 918 604 994
rect 638 918 650 994
rect 592 906 650 918
rect 850 994 908 1006
rect 850 918 862 994
rect 896 918 908 994
rect 850 906 908 918
rect 1008 918 1020 1194
rect 1054 918 1066 1194
rect 1008 906 1066 918
rect 1266 1194 1324 1206
rect 1266 918 1278 1194
rect 1312 918 1324 1194
rect 1266 906 1324 918
rect 1424 1194 1482 1206
rect 1424 918 1436 1194
rect 1470 918 1482 1194
rect 1424 906 1482 918
rect 1682 1194 1740 1206
rect 1682 918 1694 1194
rect 1728 918 1740 1194
rect 1682 906 1740 918
<< mvndiffc >>
rect 1258 2080 1292 2256
rect 1416 2080 1450 2256
rect 3472 2080 3506 2256
rect 3630 2080 3664 2256
rect 5686 2080 5720 2256
rect 5844 2080 5878 2256
rect 188 382 222 458
rect 446 382 480 458
rect 604 382 638 458
rect 862 382 896 458
rect 1020 282 1054 458
rect 1278 282 1312 458
rect 1436 282 1470 458
rect 1694 282 1728 458
<< mvpdiffc >>
rect 188 918 222 994
rect 446 918 480 994
rect 604 918 638 994
rect 862 918 896 994
rect 1020 918 1054 1194
rect 1278 918 1312 1194
rect 1436 918 1470 1194
rect 1694 918 1728 1194
<< mvpsubdiff >>
rect 2026 2918 2050 2952
rect 6336 2918 6488 2952
rect 1110 2478 1598 2490
rect 1110 2444 1218 2478
rect 1490 2444 1598 2478
rect 1110 2432 1598 2444
rect 1110 2382 1168 2432
rect 1110 1954 1122 2382
rect 1156 1954 1168 2382
rect 1540 2382 1598 2432
rect 1110 1904 1168 1954
rect 1540 1954 1552 2382
rect 1586 1954 1598 2382
rect 1540 1904 1598 1954
rect 1110 1892 1598 1904
rect 1110 1858 1218 1892
rect 1490 1858 1598 1892
rect 1110 1846 1598 1858
rect 3324 2478 3812 2490
rect 3324 2444 3432 2478
rect 3704 2444 3812 2478
rect 3324 2432 3812 2444
rect 3324 2382 3382 2432
rect 3324 1954 3336 2382
rect 3370 1954 3382 2382
rect 3754 2382 3812 2432
rect 3324 1904 3382 1954
rect 3754 1954 3766 2382
rect 3800 1954 3812 2382
rect 3754 1904 3812 1954
rect 3324 1892 3812 1904
rect 3324 1858 3432 1892
rect 3704 1858 3812 1892
rect 3324 1846 3812 1858
rect 5538 2478 6026 2490
rect 5538 2444 5646 2478
rect 5918 2444 6026 2478
rect 5538 2432 6026 2444
rect 5538 2382 5596 2432
rect 5538 1954 5550 2382
rect 5584 1954 5596 2382
rect 5968 2382 6026 2432
rect 5538 1904 5596 1954
rect 5968 1954 5980 2382
rect 6014 1954 6026 2382
rect 5968 1904 6026 1954
rect 5538 1892 6026 1904
rect 5538 1858 5646 1892
rect 5918 1858 6026 1892
rect 5538 1846 6026 1858
rect 2026 1384 2050 1418
rect 6336 1384 6488 1418
rect 42 584 100 608
rect 42 156 54 584
rect 88 156 100 584
rect 1816 584 1874 608
rect 42 106 100 156
rect 1816 156 1828 584
rect 1862 156 1874 584
rect 1816 106 1874 156
rect 42 94 1874 106
rect 42 60 148 94
rect 1768 60 1874 94
rect 42 48 1874 60
<< mvnsubdiff >>
rect 834 2746 1874 2766
rect 834 2712 916 2746
rect 1792 2712 1874 2746
rect 834 2691 1874 2712
rect 834 2684 910 2691
rect 834 1652 854 2684
rect 888 1652 910 2684
rect 1798 2684 1874 2691
rect 834 1645 910 1652
rect 1798 1652 1820 2684
rect 1854 1652 1874 2684
rect 1798 1645 1874 1652
rect 834 1624 1874 1645
rect 834 1590 916 1624
rect 1792 1590 1874 1624
rect 834 1570 1874 1590
rect 3048 2746 4088 2766
rect 3048 2712 3130 2746
rect 4006 2712 4088 2746
rect 3048 2692 4088 2712
rect 3048 2686 3122 2692
rect 3048 1650 3068 2686
rect 3102 1650 3122 2686
rect 4013 2686 4088 2692
rect 3048 1644 3122 1650
rect 4013 1650 4034 2686
rect 4068 1650 4088 2686
rect 4013 1644 4088 1650
rect 3048 1624 4088 1644
rect 3048 1590 3130 1624
rect 4006 1590 4088 1624
rect 3048 1570 4088 1590
rect 5262 2746 6302 2766
rect 5262 2712 5344 2746
rect 6220 2712 6302 2746
rect 5262 2692 6302 2712
rect 5262 2686 5336 2692
rect 5262 1650 5282 2686
rect 5316 1650 5336 2686
rect 6228 2686 6302 2692
rect 5262 1644 5336 1650
rect 6228 1650 6248 2686
rect 6282 1650 6302 2686
rect 6228 1644 6302 1650
rect 5262 1624 6302 1644
rect 5262 1590 5344 1624
rect 6220 1590 6302 1624
rect 5262 1570 6302 1590
rect 42 1426 1874 1438
rect 42 1392 148 1426
rect 1766 1392 1874 1426
rect 42 1380 1874 1392
rect 42 1330 100 1380
rect 42 784 54 1330
rect 88 784 100 1330
rect 1816 1330 1874 1380
rect 42 760 100 784
rect 1816 784 1828 1330
rect 1862 784 1874 1330
rect 1816 760 1874 784
<< mvpsubdiffcont >>
rect 2050 2918 6336 2952
rect 1218 2444 1490 2478
rect 1122 1954 1156 2382
rect 1552 1954 1586 2382
rect 1218 1858 1490 1892
rect 3432 2444 3704 2478
rect 3336 1954 3370 2382
rect 3766 1954 3800 2382
rect 3432 1858 3704 1892
rect 5646 2444 5918 2478
rect 5550 1954 5584 2382
rect 5980 1954 6014 2382
rect 5646 1858 5918 1892
rect 6454 1418 6488 2918
rect 2050 1384 6336 1418
rect 54 156 88 584
rect 1828 156 1862 584
rect 148 60 1768 94
<< mvnsubdiffcont >>
rect 916 2712 1792 2746
rect 854 1652 888 2684
rect 1820 1652 1854 2684
rect 916 1590 1792 1624
rect 3130 2712 4006 2746
rect 3068 1650 3102 2686
rect 4034 1650 4068 2686
rect 3130 1590 4006 1624
rect 5344 2712 6220 2746
rect 5282 1650 5316 2686
rect 6248 1650 6282 2686
rect 5344 1590 6220 1624
rect 148 1392 1766 1426
rect 54 784 88 1330
rect 1828 784 1862 1330
<< poly >>
rect 1304 2340 1404 2356
rect 1304 2306 1320 2340
rect 1388 2306 1404 2340
rect 1304 2268 1404 2306
rect 1304 2030 1404 2068
rect 1304 1996 1320 2030
rect 1388 1996 1404 2030
rect 1304 1980 1404 1996
rect 3518 2340 3618 2356
rect 3518 2306 3534 2340
rect 3602 2306 3618 2340
rect 3518 2268 3618 2306
rect 3518 2030 3618 2068
rect 3518 1996 3534 2030
rect 3602 1996 3618 2030
rect 3518 1980 3618 1996
rect 5732 2340 5832 2356
rect 5732 2306 5748 2340
rect 5816 2306 5832 2340
rect 5732 2268 5832 2306
rect 5732 2030 5832 2068
rect 5732 1996 5748 2030
rect 5816 1996 5832 2030
rect 5732 1980 5832 1996
rect 1066 1288 1266 1304
rect 1066 1254 1082 1288
rect 1250 1254 1266 1288
rect 1066 1206 1266 1254
rect 1482 1288 1682 1304
rect 1482 1254 1498 1288
rect 1666 1254 1682 1288
rect 1482 1206 1682 1254
rect 234 1088 434 1104
rect 234 1054 250 1088
rect 418 1054 434 1088
rect 234 1006 434 1054
rect 650 1088 850 1104
rect 650 1054 666 1088
rect 834 1054 850 1088
rect 650 1006 850 1054
rect 234 858 434 906
rect 234 824 250 858
rect 418 824 434 858
rect 234 808 434 824
rect 650 858 850 906
rect 650 824 666 858
rect 834 824 850 858
rect 650 808 850 824
rect 1066 858 1266 906
rect 1066 824 1082 858
rect 1250 824 1266 858
rect 1066 808 1266 824
rect 1482 858 1682 906
rect 1482 824 1498 858
rect 1666 824 1682 858
rect 1482 808 1682 824
rect 234 542 434 558
rect 234 508 250 542
rect 418 508 434 542
rect 234 470 434 508
rect 650 542 850 558
rect 650 508 666 542
rect 834 508 850 542
rect 650 470 850 508
rect 1066 542 1266 558
rect 1066 508 1082 542
rect 1250 508 1266 542
rect 1066 470 1266 508
rect 1482 542 1682 558
rect 1482 508 1498 542
rect 1666 508 1682 542
rect 1482 470 1682 508
rect 234 332 434 370
rect 234 298 250 332
rect 418 298 434 332
rect 234 282 434 298
rect 650 332 850 370
rect 650 298 666 332
rect 834 298 850 332
rect 650 282 850 298
rect 1066 232 1266 270
rect 1066 198 1082 232
rect 1250 198 1266 232
rect 1066 182 1266 198
rect 1482 232 1682 270
rect 1482 198 1498 232
rect 1666 198 1682 232
rect 1482 182 1682 198
<< polycont >>
rect 1320 2306 1388 2340
rect 1320 1996 1388 2030
rect 3534 2306 3602 2340
rect 3534 1996 3602 2030
rect 5748 2306 5816 2340
rect 5748 1996 5816 2030
rect 1082 1254 1250 1288
rect 1498 1254 1666 1288
rect 250 1054 418 1088
rect 666 1054 834 1088
rect 250 824 418 858
rect 666 824 834 858
rect 1082 824 1250 858
rect 1498 824 1666 858
rect 250 508 418 542
rect 666 508 834 542
rect 1082 508 1250 542
rect 1498 508 1666 542
rect 250 298 418 332
rect 666 298 834 332
rect 1082 198 1250 232
rect 1498 198 1666 232
<< locali >>
rect 2034 2918 2050 2952
rect 6336 2918 6488 2952
rect 854 2712 916 2746
rect 1792 2712 1854 2746
rect 854 2684 888 2712
rect 1820 2684 1854 2712
rect 1122 2444 1218 2478
rect 1490 2444 1586 2478
rect 1122 2382 1156 2444
rect 1552 2382 1586 2444
rect 1304 2306 1320 2340
rect 1388 2306 1404 2340
rect 1258 2256 1292 2272
rect 1258 2064 1292 2080
rect 1416 2256 1450 2272
rect 1416 2064 1450 2080
rect 1304 1996 1320 2030
rect 1388 1996 1404 2030
rect 1122 1892 1156 1954
rect 1552 1892 1586 1954
rect 1122 1858 1218 1892
rect 1490 1858 1586 1892
rect 854 1624 888 1652
rect 1820 1624 1854 1652
rect 854 1590 916 1624
rect 1792 1590 1854 1624
rect 3068 2712 3130 2746
rect 4006 2712 4068 2746
rect 3068 2686 3102 2712
rect 4034 2686 4068 2712
rect 3336 2444 3432 2478
rect 3704 2444 3800 2478
rect 3336 2382 3370 2444
rect 3766 2382 3800 2444
rect 3518 2306 3534 2340
rect 3602 2306 3618 2340
rect 3472 2256 3506 2272
rect 3472 2064 3506 2080
rect 3630 2256 3664 2272
rect 3630 2064 3664 2080
rect 3518 1996 3534 2030
rect 3602 1996 3618 2030
rect 3336 1892 3370 1954
rect 3766 1892 3800 1954
rect 3336 1858 3432 1892
rect 3704 1858 3800 1892
rect 3068 1624 3102 1650
rect 4034 1624 4068 1650
rect 3068 1590 3130 1624
rect 4006 1590 4068 1624
rect 5282 2712 5344 2746
rect 6220 2712 6282 2746
rect 5282 2686 5316 2712
rect 6248 2686 6282 2712
rect 5550 2444 5646 2478
rect 5918 2444 6014 2478
rect 5550 2382 5584 2444
rect 5980 2382 6014 2444
rect 5732 2306 5748 2340
rect 5816 2306 5832 2340
rect 5686 2256 5720 2272
rect 5686 2064 5720 2080
rect 5844 2256 5878 2272
rect 5844 2064 5878 2080
rect 5732 1996 5748 2030
rect 5816 1996 5832 2030
rect 5550 1892 5584 1954
rect 5980 1892 6014 1954
rect 5550 1858 5646 1892
rect 5918 1858 6014 1892
rect 5282 1624 5316 1650
rect 6248 1624 6282 1650
rect 5282 1590 5344 1624
rect 6220 1590 6282 1624
rect 54 1392 148 1426
rect 1766 1392 1862 1426
rect 54 1330 88 1392
rect 1828 1330 1862 1392
rect 2034 1384 2050 1418
rect 6336 1384 6488 1418
rect 1066 1254 1082 1288
rect 1250 1254 1266 1288
rect 1482 1254 1498 1288
rect 1666 1254 1682 1288
rect 1020 1194 1054 1210
rect 234 1054 250 1088
rect 418 1054 434 1088
rect 650 1054 666 1088
rect 834 1054 850 1088
rect 188 994 222 1010
rect 188 902 222 918
rect 446 994 480 1010
rect 446 902 480 918
rect 604 994 638 1010
rect 604 902 638 918
rect 862 994 986 1010
rect 896 918 986 994
rect 862 902 986 918
rect 1020 902 1054 918
rect 1278 1194 1312 1210
rect 1278 902 1312 918
rect 1436 1194 1470 1210
rect 1436 902 1470 918
rect 1694 1194 1728 1210
rect 1694 902 1728 918
rect 896 858 986 902
rect 234 824 250 858
rect 418 824 434 858
rect 650 824 666 858
rect 834 824 850 858
rect 896 824 1082 858
rect 1250 824 1266 858
rect 1482 824 1498 858
rect 1666 824 1682 858
rect 54 768 88 784
rect 54 584 88 600
rect 896 542 1266 824
rect 1828 768 1862 784
rect 1828 584 1862 600
rect 234 508 250 542
rect 418 508 434 542
rect 650 508 666 542
rect 834 508 850 542
rect 896 508 1082 542
rect 1250 508 1266 542
rect 1482 508 1498 542
rect 1666 508 1682 542
rect 896 474 986 508
rect 188 458 222 474
rect 188 366 222 382
rect 446 458 480 474
rect 446 366 480 382
rect 604 458 638 474
rect 604 366 638 382
rect 862 458 986 474
rect 896 382 986 458
rect 862 366 986 382
rect 1020 458 1054 474
rect 234 298 250 332
rect 418 298 434 332
rect 650 298 666 332
rect 834 298 850 332
rect 1020 266 1054 282
rect 1278 458 1312 474
rect 1278 266 1312 282
rect 1436 458 1470 474
rect 1436 266 1470 282
rect 1694 458 1728 474
rect 1694 266 1728 282
rect 1066 198 1082 232
rect 1250 198 1266 232
rect 1482 198 1498 232
rect 1666 198 1682 232
rect 54 94 88 156
rect 1828 94 1862 156
rect 54 60 148 94
rect 1768 60 1862 94
<< viali >>
rect 2050 2918 6336 2952
rect 942 2712 1766 2746
rect 854 1652 888 2684
rect 1218 2444 1490 2478
rect 1122 2312 1156 2382
rect 1320 2306 1388 2340
rect 1258 2080 1292 2256
rect 1416 2080 1450 2256
rect 1122 1954 1156 2024
rect 1320 1996 1388 2030
rect 1552 1954 1586 2382
rect 1218 1858 1490 1892
rect 1820 1652 1854 2684
rect 942 1590 1766 1624
rect 3156 2712 3980 2746
rect 3068 1652 3102 2684
rect 3432 2444 3704 2478
rect 3336 2312 3370 2382
rect 3534 2306 3602 2340
rect 3472 2080 3506 2256
rect 3630 2080 3664 2256
rect 3336 1954 3370 2024
rect 3534 1996 3602 2030
rect 3766 1954 3800 2382
rect 3432 1858 3704 1892
rect 4034 1652 4068 2684
rect 3156 1590 3980 1624
rect 5370 2712 6194 2746
rect 5282 1652 5316 2684
rect 5646 2444 5918 2478
rect 5550 2312 5584 2382
rect 5748 2306 5816 2340
rect 5686 2080 5720 2256
rect 5844 2080 5878 2256
rect 5550 1954 5584 2024
rect 5748 1996 5816 2030
rect 5980 1954 6014 2382
rect 5646 1858 5918 1892
rect 6248 1652 6282 2684
rect 5370 1590 6194 1624
rect 148 1392 1766 1426
rect 6454 1418 6488 2918
rect 54 784 88 1330
rect 2050 1384 6336 1418
rect 1082 1254 1250 1288
rect 1498 1254 1666 1288
rect 250 1054 418 1088
rect 666 1054 834 1088
rect 188 918 222 994
rect 446 918 480 994
rect 604 918 638 994
rect 862 918 896 994
rect 1020 918 1054 1194
rect 1278 918 1312 1194
rect 1436 918 1470 1194
rect 1694 918 1728 1194
rect 250 824 418 858
rect 666 824 834 858
rect 1082 824 1250 858
rect 1498 824 1666 858
rect 54 156 88 584
rect 1828 784 1862 1330
rect 250 508 418 542
rect 666 508 834 542
rect 1082 508 1250 542
rect 1498 508 1666 542
rect 188 382 222 458
rect 446 382 480 458
rect 604 382 638 458
rect 862 382 896 458
rect 250 298 418 332
rect 666 298 834 332
rect 1020 282 1054 458
rect 1278 282 1312 458
rect 1436 282 1470 458
rect 1694 282 1728 458
rect 1082 198 1250 232
rect 1498 198 1666 232
rect 1828 156 1862 584
rect 148 60 1768 94
<< metal1 >>
rect 2038 2952 6494 2958
rect 2038 2918 2050 2952
rect 6336 2918 6494 2952
rect 2038 2912 6454 2918
rect 848 2746 1860 2752
rect 848 2712 942 2746
rect 1766 2712 1860 2746
rect 848 2706 1860 2712
rect 848 2684 894 2706
rect 848 1652 854 2684
rect 888 1652 894 2684
rect 1814 2684 1860 2706
rect 1116 2478 1592 2484
rect 1116 2444 1218 2478
rect 1490 2444 1592 2478
rect 1116 2382 1592 2444
rect 1116 2312 1122 2382
rect 1156 2340 1552 2382
rect 1156 2312 1320 2340
rect 1116 2306 1320 2312
rect 1388 2306 1552 2340
rect 1116 2300 1552 2306
rect 1116 2256 1298 2268
rect 1292 2080 1298 2256
rect 1116 2068 1298 2080
rect 1410 2256 1552 2300
rect 1586 2256 1592 2382
rect 1410 2080 1416 2256
rect 1410 2036 1552 2080
rect 1116 2030 1552 2036
rect 1116 2024 1320 2030
rect 1116 1954 1122 2024
rect 1156 1996 1320 2024
rect 1388 1996 1552 2030
rect 1156 1954 1552 1996
rect 1586 1954 1592 2080
rect 1116 1892 1592 1954
rect 1116 1858 1218 1892
rect 1490 1858 1592 1892
rect 1116 1852 1592 1858
rect 1814 1736 1820 2684
rect 848 1630 894 1652
rect 1660 1730 1820 1736
rect 1660 1630 1666 1730
rect 848 1624 1666 1630
rect 848 1590 942 1624
rect 848 1584 1666 1590
rect 48 1542 1666 1584
rect 1854 1542 1860 2684
rect 48 1432 1860 1542
rect 3062 2746 4074 2752
rect 3062 2712 3156 2746
rect 3980 2712 4074 2746
rect 3062 2706 4074 2712
rect 3062 2684 3108 2706
rect 3062 1542 3068 2684
rect 3102 1736 3108 2684
rect 4028 2684 4074 2706
rect 3330 2478 3806 2484
rect 3330 2444 3432 2478
rect 3704 2444 3806 2478
rect 3330 2382 3806 2444
rect 3330 2312 3336 2382
rect 3370 2340 3766 2382
rect 3370 2312 3534 2340
rect 3330 2306 3534 2312
rect 3602 2306 3766 2340
rect 3330 2300 3766 2306
rect 3330 2256 3512 2268
rect 3506 2080 3512 2256
rect 3330 2068 3512 2080
rect 3624 2256 3766 2300
rect 3800 2256 3806 2382
rect 3624 2080 3630 2256
rect 3624 2036 3766 2080
rect 3330 2030 3766 2036
rect 3330 2024 3534 2030
rect 3330 1954 3336 2024
rect 3370 1996 3534 2024
rect 3602 1996 3766 2030
rect 3370 1954 3766 1996
rect 3800 1954 3806 2080
rect 3330 1892 3806 1954
rect 3330 1858 3432 1892
rect 3704 1858 3806 1892
rect 3330 1852 3806 1858
rect 3102 1730 3262 1736
rect 3256 1630 3262 1730
rect 4028 1652 4034 2684
rect 4068 1652 4074 2684
rect 4028 1630 4074 1652
rect 3256 1624 4074 1630
rect 3980 1590 4074 1624
rect 3256 1584 4074 1590
rect 5276 2746 6288 2752
rect 5276 2712 5370 2746
rect 6194 2712 6288 2746
rect 5276 2706 6288 2712
rect 5276 2684 5322 2706
rect 3256 1542 3262 1584
rect 3062 1536 3262 1542
rect 5276 1542 5282 2684
rect 5316 1736 5322 2684
rect 6242 2684 6288 2706
rect 5544 2478 6020 2484
rect 5544 2444 5646 2478
rect 5918 2444 6020 2478
rect 5544 2382 6020 2444
rect 5544 2312 5550 2382
rect 5584 2340 5980 2382
rect 5584 2312 5748 2340
rect 5544 2306 5748 2312
rect 5816 2306 5980 2340
rect 5544 2300 5980 2306
rect 5544 2256 5726 2268
rect 5720 2080 5726 2256
rect 5544 2068 5726 2080
rect 5838 2256 5980 2300
rect 6014 2256 6020 2382
rect 5838 2080 5844 2256
rect 5838 2036 5980 2080
rect 5544 2030 5980 2036
rect 5544 2024 5748 2030
rect 5544 1954 5550 2024
rect 5584 1996 5748 2024
rect 5816 1996 5980 2030
rect 5584 1954 5980 1996
rect 6014 1954 6020 2080
rect 5544 1892 6020 1954
rect 5544 1858 5646 1892
rect 5918 1858 6020 1892
rect 5544 1852 6020 1858
rect 5316 1730 5476 1736
rect 5470 1630 5476 1730
rect 6242 1652 6248 2684
rect 6282 1652 6288 2684
rect 6242 1630 6288 1652
rect 5470 1624 6288 1630
rect 6194 1590 6288 1624
rect 5470 1584 6288 1590
rect 5470 1542 5476 1584
rect 5276 1536 5476 1542
rect 48 1426 1868 1432
rect 6448 1426 6454 2912
rect 48 1392 148 1426
rect 1766 1392 1868 1426
rect 48 1386 1868 1392
rect 48 1330 1048 1386
rect 48 784 54 1330
rect 88 1218 1048 1330
rect 1076 1288 1256 1300
rect 1076 1254 1082 1288
rect 1250 1254 1256 1288
rect 1076 1242 1256 1254
rect 88 1194 1060 1218
rect 88 1128 1020 1194
rect 88 1006 216 1128
rect 244 1088 424 1100
rect 244 1054 250 1088
rect 418 1054 424 1088
rect 244 1042 424 1054
rect 88 994 228 1006
rect 88 918 188 994
rect 222 918 228 994
rect 88 906 228 918
rect 88 784 94 906
rect 256 870 412 1042
rect 564 1018 632 1128
rect 660 1088 840 1100
rect 660 1054 666 1088
rect 834 1054 840 1088
rect 660 1042 840 1054
rect 440 994 536 1006
rect 440 918 446 994
rect 480 918 536 994
rect 440 906 536 918
rect 564 994 644 1018
rect 564 918 604 994
rect 638 918 644 994
rect 564 906 644 918
rect 48 772 94 784
rect 244 858 424 870
rect 244 824 250 858
rect 418 824 424 858
rect 244 734 424 824
rect 48 634 424 734
rect 48 584 94 596
rect 48 248 54 584
rect 42 242 54 248
rect 88 470 94 584
rect 244 542 424 634
rect 244 508 250 542
rect 418 508 424 542
rect 244 496 424 508
rect 486 772 536 906
rect 672 870 828 1042
rect 856 994 902 1006
rect 856 918 862 994
rect 896 918 902 994
rect 856 906 902 918
rect 930 918 1020 1128
rect 1054 918 1060 1194
rect 930 906 1060 918
rect 1088 870 1244 1242
rect 1358 1210 1464 1386
rect 1822 1330 1868 1386
rect 2038 1374 2050 1426
rect 6488 1418 6494 2918
rect 6466 1374 6494 1418
rect 1492 1288 1672 1300
rect 1492 1254 1498 1288
rect 1666 1254 1672 1288
rect 1492 1242 1672 1254
rect 1272 1194 1330 1206
rect 1272 918 1278 1194
rect 1272 906 1330 918
rect 1358 1194 1476 1210
rect 1358 918 1436 1194
rect 1470 918 1476 1194
rect 1358 906 1476 918
rect 1504 870 1660 1242
rect 1688 1194 1746 1206
rect 1688 918 1694 1194
rect 1688 906 1746 918
rect 660 858 840 870
rect 660 824 666 858
rect 834 824 840 858
rect 660 772 840 824
rect 1076 858 1256 870
rect 1076 824 1082 858
rect 1250 824 1256 858
rect 1076 812 1256 824
rect 1492 858 1672 870
rect 1492 824 1498 858
rect 1666 824 1672 858
rect 1492 772 1672 824
rect 1822 784 1828 1330
rect 1862 784 1868 1330
rect 1822 772 1868 784
rect 486 594 1672 772
rect 88 458 228 470
rect 88 382 188 458
rect 222 382 228 458
rect 88 370 228 382
rect 88 258 216 370
rect 256 344 412 496
rect 486 470 536 594
rect 660 542 840 594
rect 660 508 666 542
rect 834 508 840 542
rect 660 496 840 508
rect 1076 542 1256 554
rect 1076 508 1082 542
rect 1250 508 1256 542
rect 1076 496 1256 508
rect 1492 542 1672 594
rect 1492 508 1498 542
rect 1666 508 1672 542
rect 1492 496 1672 508
rect 1822 584 1868 596
rect 440 458 536 470
rect 440 382 446 458
rect 480 382 536 458
rect 440 370 536 382
rect 564 458 644 470
rect 564 382 604 458
rect 638 382 644 458
rect 564 368 644 382
rect 244 332 424 344
rect 244 298 250 332
rect 418 298 424 332
rect 244 286 424 298
rect 564 258 632 368
rect 672 344 828 496
rect 856 458 902 470
rect 856 382 862 458
rect 896 382 902 458
rect 856 370 902 382
rect 930 458 1060 470
rect 660 332 840 344
rect 660 298 666 332
rect 834 298 840 332
rect 660 286 840 298
rect 930 282 1020 458
rect 1054 282 1060 458
rect 930 268 1060 282
rect 930 258 1048 268
rect 88 242 1048 258
rect 1088 244 1244 496
rect 1272 458 1330 470
rect 1272 282 1278 458
rect 1272 270 1330 282
rect 1358 458 1476 470
rect 1358 282 1436 458
rect 1470 282 1476 458
rect 1358 270 1476 282
rect 42 54 48 242
rect 236 100 1048 242
rect 1076 232 1256 244
rect 1076 198 1082 232
rect 1250 198 1256 232
rect 1076 186 1256 198
rect 1358 100 1464 270
rect 1504 244 1660 496
rect 1688 458 1746 470
rect 1688 282 1694 458
rect 1688 270 1746 282
rect 1492 232 1672 244
rect 1492 198 1498 232
rect 1666 198 1672 232
rect 1492 186 1672 198
rect 1822 156 1828 584
rect 1862 156 1868 584
rect 1822 100 1868 156
rect 236 94 1868 100
rect 1768 60 1868 94
rect 236 54 1868 60
rect 42 48 242 54
<< via1 >>
rect 1116 2080 1258 2256
rect 1258 2080 1292 2256
rect 1416 2080 1450 2256
rect 1450 2080 1552 2256
rect 1552 2080 1586 2256
rect 1586 2080 1592 2256
rect 1666 1652 1820 1730
rect 1820 1652 1854 1730
rect 1666 1624 1854 1652
rect 1666 1590 1766 1624
rect 1766 1590 1854 1624
rect 1666 1542 1854 1590
rect 3330 2080 3472 2256
rect 3472 2080 3506 2256
rect 3630 2080 3664 2256
rect 3664 2080 3766 2256
rect 3766 2080 3800 2256
rect 3800 2080 3806 2256
rect 3068 1652 3102 1730
rect 3102 1652 3256 1730
rect 3068 1624 3256 1652
rect 3068 1590 3156 1624
rect 3156 1590 3256 1624
rect 3068 1542 3256 1590
rect 5544 2080 5686 2256
rect 5686 2080 5720 2256
rect 5844 2080 5878 2256
rect 5878 2080 5980 2256
rect 5980 2080 6014 2256
rect 6014 2080 6020 2256
rect 5282 1652 5316 1730
rect 5316 1652 5470 1730
rect 5282 1624 5470 1652
rect 5282 1590 5370 1624
rect 5370 1590 5470 1624
rect 5282 1542 5470 1590
rect 2050 1418 6454 1426
rect 6454 1418 6466 1426
rect 2050 1384 6336 1418
rect 6336 1384 6466 1418
rect 2050 1374 6466 1384
rect 1278 918 1312 1194
rect 1312 918 1330 1194
rect 1694 918 1728 1194
rect 1728 918 1746 1194
rect 1278 282 1312 458
rect 1312 282 1330 458
rect 48 156 54 242
rect 54 156 88 242
rect 88 156 236 242
rect 48 94 236 156
rect 1694 282 1728 458
rect 1728 282 1746 458
rect 48 60 148 94
rect 148 60 236 94
rect 48 54 236 60
<< metal2 >>
rect 564 4442 764 4452
rect 564 4378 574 4442
rect 754 4378 764 4442
rect 564 3084 764 4378
rect 4596 4442 4796 4452
rect 4596 4378 4606 4442
rect 4786 4378 4796 4442
rect 564 2884 1610 3084
rect 1410 2262 1610 2884
rect 4596 2262 4796 4378
rect 1098 2256 1298 2262
rect 1098 2080 1116 2256
rect 1292 2080 1298 2256
rect 1098 1480 1298 2080
rect 1410 2256 3512 2262
rect 1410 2080 1416 2256
rect 1592 2080 3330 2256
rect 3506 2080 3512 2256
rect 1410 2074 3512 2080
rect 3624 2256 5726 2262
rect 3624 2080 3630 2256
rect 3806 2080 5544 2256
rect 5720 2080 5726 2256
rect 3624 2074 5726 2080
rect 5838 2256 6408 2262
rect 5838 2080 5844 2256
rect 6020 2080 6408 2256
rect 5838 2074 6408 2080
rect 6472 2074 6482 2262
rect 1660 1730 5476 1736
rect 1660 1542 1666 1730
rect 1854 1542 3068 1730
rect 3256 1542 5282 1730
rect 5470 1542 5476 1730
rect 1660 1536 5476 1542
rect 720 1474 6482 1480
rect 720 1426 6408 1474
rect 720 1374 2050 1426
rect 720 1286 6408 1374
rect 6472 1286 6482 1474
rect 720 1280 6482 1286
rect 720 248 920 1280
rect 42 242 920 248
rect 42 54 48 242
rect 236 54 920 242
rect 42 48 920 54
rect 1272 1194 1336 1200
rect 1272 918 1278 1194
rect 1330 918 1336 1194
rect 1272 470 1336 918
rect 1688 1194 1752 1200
rect 1688 918 1694 1194
rect 1746 918 1752 1194
rect 1688 470 1752 918
rect 1272 458 1472 470
rect 1272 282 1278 458
rect 1330 282 1472 458
rect 1272 -924 1472 282
rect 496 -1124 1472 -924
rect 1688 458 1888 470
rect 1688 282 1694 458
rect 1746 282 1888 458
rect 496 -1408 696 -1124
rect 496 -1472 506 -1408
rect 686 -1472 696 -1408
rect 496 -1482 696 -1472
rect 1688 -1408 1888 282
rect 1688 -1472 1698 -1408
rect 1878 -1472 1888 -1408
rect 1688 -1482 1888 -1472
<< via2 >>
rect 574 4378 754 4442
rect 4606 4378 4786 4442
rect 6408 2074 6472 2262
rect 6408 1426 6472 1474
rect 6408 1374 6466 1426
rect 6466 1374 6472 1426
rect 6408 1286 6472 1374
rect 506 -1472 686 -1408
rect 1698 -1472 1878 -1408
<< metal3 >>
rect 568 4442 770 4448
rect 4600 4442 4796 4448
rect -4266 4378 -4260 4442
rect 764 4378 770 4442
rect 1074 4378 1080 4442
rect 6104 4378 6110 4442
rect 568 4372 770 4378
rect 4600 4372 4796 4378
rect -4288 4272 792 4292
rect -4288 4208 -4260 4272
rect 764 4208 792 4272
rect -4288 -1140 792 4208
rect 1052 4272 6132 4292
rect 1052 4208 1080 4272
rect 6104 4208 6132 4272
rect 1052 -1140 6132 4208
rect 6408 3854 6472 3860
rect 6402 2068 6408 2268
rect 6472 2068 6478 2268
rect 6408 1614 6472 1620
rect 6408 1528 6472 1534
rect 6402 1280 6408 1480
rect 6558 1528 12990 3940
rect 6472 1280 6478 1480
rect 6408 -1118 6472 -1112
rect 6558 -1112 6578 1528
rect 6642 -1112 12990 1528
rect 6558 -1140 12990 -1112
rect 496 -1408 702 -1402
rect 1692 -1408 1884 -1402
rect -4198 -1472 -4192 -1408
rect 696 -1472 702 -1408
rect 1142 -1472 1148 -1408
rect 6036 -1472 6042 -1408
rect 496 -1478 702 -1472
rect 1692 -1478 1884 -1472
<< via3 >>
rect -4260 4378 574 4442
rect 574 4378 754 4442
rect 754 4378 764 4442
rect 1080 4378 4606 4442
rect 4606 4378 4786 4442
rect 4786 4378 6104 4442
rect -4260 4208 764 4272
rect 1080 4208 6104 4272
rect 6408 2262 6472 3854
rect 6408 2074 6472 2262
rect 6408 1620 6472 2074
rect 6408 1474 6472 1528
rect 6408 1286 6472 1474
rect 6408 -1112 6472 1286
rect 6578 -1112 6642 1528
rect -4192 -1472 506 -1408
rect 506 -1472 686 -1408
rect 686 -1472 696 -1408
rect 1148 -1472 1698 -1408
rect 1698 -1472 1878 -1408
rect 1878 -1472 6036 -1408
<< mimcap >>
rect -4248 3860 752 3900
rect -4248 -1060 -4208 3860
rect 712 -1060 752 3860
rect -4248 -1100 752 -1060
rect 1092 3860 6092 3900
rect 1092 -1060 1132 3860
rect 6052 -1060 6092 3860
rect 1092 -1100 6092 -1060
rect 6950 3860 12950 3900
rect 6950 -1060 6990 3860
rect 12910 -1060 12950 3860
rect 6950 -1100 12950 -1060
<< mimcapcontact >>
rect -4208 -1060 712 3860
rect 1132 -1060 6052 3860
rect 6990 -1060 12910 3860
<< metal4 >>
rect -4276 4442 780 4458
rect -4276 4378 -4260 4442
rect 764 4378 780 4442
rect -4276 4272 780 4378
rect -4276 4208 -4260 4272
rect 764 4208 780 4272
rect -4276 4192 780 4208
rect 1064 4442 6120 4458
rect 1064 4378 1080 4442
rect 6104 4378 6120 4442
rect 1064 4272 6120 4378
rect 1064 4208 1080 4272
rect 6104 4208 6120 4272
rect 1064 4192 6120 4208
rect -4209 3860 713 3861
rect -4209 -1060 -4208 3860
rect 712 -1060 713 3860
rect -4209 -1061 713 -1060
rect 1131 3860 6053 3861
rect 6989 3860 12911 3861
rect 1131 -1060 1132 3860
rect 6052 -1060 6053 3860
rect 6392 3854 6990 3860
rect 6392 1620 6408 3854
rect 6472 1620 6990 3854
rect 6392 1614 6990 1620
rect 1131 -1061 6053 -1060
rect 6392 1528 6658 1534
rect -4208 -1408 712 -1061
rect -4208 -1472 -4192 -1408
rect 696 -1472 712 -1408
rect -4208 -1488 712 -1472
rect 1132 -1408 6052 -1061
rect 6392 -1112 6408 1528
rect 6472 -1112 6578 1528
rect 6642 -1112 6658 1528
rect 6989 -1060 6990 1614
rect 12910 -1060 12911 3860
rect 6989 -1061 12911 -1060
rect 6392 -1128 6658 -1112
rect 1132 -1472 1148 -1408
rect 6036 -1472 6052 -1408
rect 1132 -1488 6052 -1472
<< labels >>
flabel metal1 486 370 536 1006 0 FreeMono 160 90 0 0 clkinb
flabel locali 902 370 952 1006 0 FreeMono 160 90 0 0 clkina
flabel viali 148 1392 182 1426 0 FreeMono 160 0 0 0 VAPWR
flabel viali 1278 282 1312 458 0 FreeMono 160 90 0 0 clka
flabel viali 1278 918 1312 1194 0 FreeMono 160 90 0 0 clka
flabel viali 1694 918 1728 1194 0 FreeMono 160 90 0 0 clkb
flabel viali 1694 282 1728 458 0 FreeMono 160 90 0 0 clkb
flabel viali 1416 2080 1450 2256 0 FreeMono 160 90 0 0 stage1
flabel viali 3472 2080 3506 2256 0 FreeMono 160 90 0 0 stage1
flabel viali 3630 2080 3664 2256 0 FreeMono 160 90 0 0 stage2
flabel viali 854 1652 888 1686 0 FreeMono 160 0 0 0 VAPWR
flabel viali 5686 2080 5720 2256 0 FreeMono 160 90 0 0 stage2
flabel viali 5844 2080 5878 2256 0 FreeMono 160 90 0 0 VOUT
flabel metal4 1132 -1060 6052 3860 0 FreeMono 1600 180 0 0 clkb
flabel metal4 -4208 -1060 712 3860 0 FreeMono 1600 180 0 0 clka
flabel metal3 1052 4192 6132 4292 0 FreeMono 480 180 0 0 stage2
flabel metal3 -4288 4192 792 4292 0 FreeMono 480 180 0 0 stage1
flabel viali 2050 1384 2084 1418 0 FreeMono 160 0 0 0 VGND
flabel viali 2050 2918 2084 2952 0 FreeMono 160 0 0 0 VGND
flabel metal1 48 634 148 734 0 FreeMono 160 0 0 0 clk
port 0 nsew
flabel metal1 48 1232 248 1432 0 FreeSans 256 0 0 0 VAPWR
port 2 nsew
flabel via1 48 54 236 242 0 FreeMono 160 0 0 0 VGND
port 3 nsew
flabel viali 248 60 282 94 0 FreeMono 160 0 0 0 VGND
flabel metal4 6990 -1060 12910 3860 0 FreeMono 1600 180 0 0 VOUT
flabel metal3 6558 -1140 6578 3940 0 FreeMono 480 90 0 0 VGND
flabel metal2 6402 2074 6482 2262 0 FreeMono 320 90 0 0 VOUT
port 1 nsew
flabel viali 1320 1996 1388 2030 0 FreeMono 96 0 0 0 stage1
flabel viali 1320 2306 1388 2340 0 FreeMono 96 0 0 0 stage1
flabel viali 1258 2080 1292 2256 0 FreeMono 160 90 0 0 VGND
flabel viali 3336 1954 3370 1988 0 FreeMono 160 0 0 0 stage2
flabel viali 5550 1954 5584 1988 0 FreeMono 160 0 0 0 VOUT
flabel viali 1122 1954 1156 1988 0 FreeMono 160 0 0 0 stage1
flabel mvnsubdiffcont 3068 1650 3102 1684 0 FreeMono 160 0 0 0 VAPWR
flabel mvnsubdiffcont 5282 1650 5316 1684 0 FreeMono 160 0 0 0 VAPWR
flabel viali 3534 1996 3602 2030 0 FreeMono 96 0 0 0 stage2
flabel viali 3534 2306 3602 2340 0 FreeMono 96 0 0 0 stage2
flabel viali 5748 2306 5816 2340 0 FreeMono 96 0 0 0 VOUT
flabel viali 5748 1996 5816 2030 0 FreeMono 96 0 0 0 VOUT
<< end >>
