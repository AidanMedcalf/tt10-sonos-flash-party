** sch_path: /home/amedcalf/projects/tt10-sonos-flash-party/xschem/vprog_controller.sch
.subckt vprog_controller pos_en neg_en VOUT VDPWR VGND VPRGPOS VPRGNEG VDPWR1
*.PININFO VPRGNEG:B neg_en:I VOUT:O VDPWR:B pos_en:I VGND:B VPRGPOS:B VDPWR1:B
XM1 net1 neg_en VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=6 m=1
XM2 neg_mid_b neg_en_b VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=6 m=1
XM4 neg_mid_b net1 VPRGNEG VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.5 nf=1 m=1
XM3 net1 neg_mid_b VPRGNEG VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.5 nf=1 m=1
XM7 vintn neg_mid_b VPRGNEG VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 L=3 W=1 nf=2 m=1
XM8 net2 pos_en_b VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=3 W=1.5 nf=3 m=1
XM12 net3 pos_mid_b VPRGPOS VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 L=3 W=0.5 nf=1 m=1
XM13 pos_mid_b net3 VPRGPOS VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 L=3 W=0.5 nf=1 m=1
XM14 pos_mid_b pos_en VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=3 W=2 nf=4 m=1
XM15 net3 pos_en_b VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=3 W=2 nf=4 m=1
XM16 vintp pos_mid_b VPRGPOS VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=6 m=1
XM11 VOUT neg_mid_b net2 net2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=6 m=1
XM17 VOUT VDPWR1 vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=6 m=1
XM18 VOUT VDPWR vintn VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 L=3 W=1 nf=2 m=1
XM5 neg_en_b neg_en VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1 nf=2 m=1
XM6 neg_en_b neg_en VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=3 W=1 nf=2 m=1
XM9 pos_en_b pos_en VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=3 W=1 nf=2 m=1
XM10 pos_en_b pos_en VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1 nf=2 m=1
.ends
.end
