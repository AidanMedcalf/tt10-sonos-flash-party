magic
tech sky130A
timestamp 1740658820
<< metal4 >>
rect 10740 8700 10830 8730
rect 10710 8670 10860 8700
rect 10680 8610 10890 8670
rect 10650 8550 10860 8610
rect 10620 8490 10830 8550
rect 10590 8460 10800 8490
rect 10560 8430 10800 8460
rect 10560 8400 10770 8430
rect 10530 8370 10770 8400
rect 10530 8340 10740 8370
rect 10500 8310 10740 8340
rect 10470 8250 10710 8310
rect 10440 8220 10680 8250
rect 10440 8190 10650 8220
rect 10410 8160 10650 8190
rect 10410 8130 10620 8160
rect 10380 8100 10620 8130
rect 10350 8040 10590 8100
rect 10320 7980 10560 8040
rect 10290 7950 10530 7980
rect 10260 7920 10530 7950
rect 10260 7890 10500 7920
rect 10230 7860 10500 7890
rect 10230 7830 10470 7860
rect 10950 7830 11070 7860
rect 10200 7800 10440 7830
rect 10860 7800 11070 7830
rect 10170 7770 10440 7800
rect 10740 7770 11040 7800
rect 10170 7740 10410 7770
rect 10620 7740 11010 7770
rect 10140 7710 11010 7740
rect 10110 7680 10980 7710
rect 10110 7650 10950 7680
rect 10080 7620 10920 7650
rect 8850 7590 8880 7620
rect 10050 7590 10890 7620
rect 8790 7560 8910 7590
rect 6240 7500 6270 7530
rect 8790 7500 8940 7560
rect 10020 7530 10860 7590
rect 9990 7500 10830 7530
rect 6060 7470 6420 7500
rect 8400 7470 8430 7500
rect 6000 7440 6510 7470
rect 8340 7440 8460 7470
rect 5940 7410 6570 7440
rect 8340 7410 8490 7440
rect 5910 7380 6600 7410
rect 5880 7350 6660 7380
rect 5850 7320 6210 7350
rect 6300 7320 6690 7350
rect 7920 7320 7980 7350
rect 5820 7290 6090 7320
rect 6420 7290 6720 7320
rect 7890 7290 8010 7320
rect 5790 7260 6030 7290
rect 6480 7260 6750 7290
rect 7890 7260 8040 7290
rect 5760 7230 6000 7260
rect 6540 7230 6750 7260
rect 5760 7200 5970 7230
rect 6570 7200 6780 7230
rect 7470 7200 7530 7230
rect 5730 7170 5940 7200
rect 6600 7170 6780 7200
rect 7440 7170 7560 7200
rect 5700 7110 5910 7170
rect 6180 7140 6360 7170
rect 6600 7140 6810 7170
rect 6120 7110 6420 7140
rect 6630 7110 6810 7140
rect 5700 7080 5880 7110
rect 6090 7080 6450 7110
rect 6630 7080 6840 7110
rect 7440 7080 7590 7170
rect 5670 7050 5880 7080
rect 6060 7050 6450 7080
rect 5670 6780 5850 7050
rect 6030 7020 6480 7050
rect 6660 7020 6840 7080
rect 7350 7050 7590 7080
rect 7230 7020 7590 7050
rect 6030 6990 6180 7020
rect 6330 6990 6510 7020
rect 6000 6870 6150 6990
rect 6360 6870 6510 6990
rect 6030 6840 6210 6870
rect 6330 6840 6510 6870
rect 6660 6930 6870 7020
rect 7140 6990 7590 7020
rect 7020 6960 7590 6990
rect 6930 6930 7590 6960
rect 6660 6900 7590 6930
rect 6660 6870 7290 6900
rect 6660 6840 7200 6870
rect 6030 6810 6480 6840
rect 6060 6780 6480 6810
rect 6660 6810 7110 6840
rect 6660 6780 7020 6810
rect 5670 6750 5880 6780
rect 6060 6750 6450 6780
rect 6660 6750 6870 6780
rect 5700 6720 5880 6750
rect 6090 6720 6420 6750
rect 5700 6690 5910 6720
rect 6150 6690 6390 6720
rect 6630 6690 6810 6750
rect 5730 6660 5910 6690
rect 6210 6660 6330 6690
rect 6600 6660 6810 6690
rect 5730 6630 5940 6660
rect 6600 6630 6780 6660
rect 5760 6600 5970 6630
rect 6570 6600 6780 6630
rect 5760 6570 6000 6600
rect 6510 6570 6750 6600
rect 5790 6540 6030 6570
rect 6480 6540 6720 6570
rect 5820 6510 6120 6540
rect 6420 6510 6720 6540
rect 5850 6480 6690 6510
rect 5880 6450 6660 6480
rect 5910 6420 6600 6450
rect 5940 6390 6570 6420
rect 6000 6360 6510 6390
rect 6090 6330 6420 6360
rect 6180 6180 6330 6330
rect 6180 5550 6360 6180
rect 7440 5910 7590 6900
rect 7860 6840 8040 7260
rect 7890 6570 8040 6840
rect 7860 6060 8040 6570
rect 8310 6240 8490 7410
rect 8760 7350 8940 7500
rect 9960 7470 10440 7500
rect 10500 7470 10800 7500
rect 9960 7440 10350 7470
rect 10470 7440 10770 7470
rect 9930 7410 10290 7440
rect 10440 7410 10740 7440
rect 9900 7380 10170 7410
rect 10440 7380 10710 7410
rect 9900 7350 10050 7380
rect 10410 7350 10710 7380
rect 8790 7200 8940 7350
rect 10380 7320 10680 7350
rect 10380 7290 10650 7320
rect 10350 7230 10620 7290
rect 8760 7080 8940 7200
rect 10320 7200 10590 7230
rect 12390 7200 12570 7230
rect 10320 7170 10560 7200
rect 12270 7170 12630 7200
rect 10290 7140 10560 7170
rect 12150 7140 12690 7170
rect 10260 7080 10530 7140
rect 12030 7110 12690 7140
rect 11940 7080 12720 7110
rect 8790 6480 8940 7080
rect 10230 7050 10500 7080
rect 11850 7050 12720 7080
rect 10230 7020 10470 7050
rect 11730 7020 12450 7050
rect 12480 7020 12720 7050
rect 10200 6990 10470 7020
rect 11640 6990 12300 7020
rect 10200 6960 10440 6990
rect 11550 6960 12210 6990
rect 10170 6930 10410 6960
rect 11460 6930 12120 6960
rect 10140 6900 10410 6930
rect 11370 6900 12030 6930
rect 12510 6900 12720 7020
rect 10140 6870 10380 6900
rect 11280 6870 11910 6900
rect 10110 6840 10350 6870
rect 11190 6840 11820 6870
rect 10080 6810 10350 6840
rect 11100 6810 11730 6840
rect 10080 6780 10320 6810
rect 11010 6780 11640 6810
rect 10050 6720 10290 6780
rect 10920 6750 11520 6780
rect 10800 6720 11430 6750
rect 10050 6690 10260 6720
rect 10710 6690 11340 6720
rect 10050 6660 10230 6690
rect 10620 6660 11250 6690
rect 10080 6630 10200 6660
rect 10530 6630 11160 6660
rect 10440 6600 11070 6630
rect 10350 6570 10980 6600
rect 10260 6540 10860 6570
rect 10170 6510 10770 6540
rect 10080 6480 10680 6510
rect 8760 6360 8940 6480
rect 9990 6450 10590 6480
rect 11730 6450 12000 6480
rect 9870 6420 10500 6450
rect 11670 6420 12120 6450
rect 9780 6390 10410 6420
rect 11610 6390 12150 6420
rect 9690 6360 10290 6390
rect 11580 6360 12120 6390
rect 8790 6330 8910 6360
rect 9600 6330 10200 6360
rect 11550 6330 12120 6360
rect 8820 6300 8880 6330
rect 9510 6300 10110 6330
rect 11520 6300 12090 6330
rect 9420 6270 10020 6300
rect 11490 6270 12090 6300
rect 9330 6240 9930 6270
rect 11490 6240 12060 6270
rect 8310 6210 8460 6240
rect 9240 6210 9840 6240
rect 11460 6210 11790 6240
rect 11940 6210 12060 6240
rect 8340 6180 8460 6210
rect 9120 6180 9720 6210
rect 11460 6180 11730 6210
rect 9030 6150 9630 6180
rect 11460 6150 11700 6180
rect 8970 6120 9540 6150
rect 8880 6090 9450 6120
rect 11430 6090 11700 6150
rect 8790 6060 9360 6090
rect 10590 6060 10890 6090
rect 11430 6060 11670 6090
rect 7890 6030 8010 6060
rect 8670 6030 9270 6060
rect 10500 6030 10980 6060
rect 7920 6000 7980 6030
rect 8580 6000 9180 6030
rect 10440 6000 11040 6030
rect 11430 6000 11700 6060
rect 8490 5970 9090 6000
rect 10380 5970 11100 6000
rect 11430 5970 11730 6000
rect 8370 5940 9000 5970
rect 10350 5940 11130 5970
rect 11430 5940 11790 5970
rect 8310 5910 8910 5940
rect 10290 5910 11160 5940
rect 11460 5910 11880 5940
rect 7470 5880 7560 5910
rect 8190 5880 8820 5910
rect 10260 5880 11190 5910
rect 11460 5880 12000 5910
rect 8130 5850 8730 5880
rect 10230 5850 11220 5880
rect 11490 5850 12060 5880
rect 8040 5820 8640 5850
rect 9840 5820 9870 5850
rect 10200 5820 10680 5850
rect 10830 5820 11250 5850
rect 11520 5820 12090 5850
rect 7920 5790 8550 5820
rect 9780 5790 9870 5820
rect 10170 5790 10560 5820
rect 10920 5790 11250 5820
rect 11550 5790 12120 5820
rect 7860 5760 8430 5790
rect 9720 5760 9870 5790
rect 7770 5730 8370 5760
rect 9660 5730 9870 5760
rect 10140 5760 10470 5790
rect 10950 5760 11280 5790
rect 11610 5760 12150 5790
rect 10140 5730 10440 5760
rect 11010 5730 11280 5760
rect 11670 5730 12180 5760
rect 7680 5700 8280 5730
rect 7560 5670 8160 5700
rect 7500 5640 8070 5670
rect 7380 5610 7980 5640
rect 7290 5580 7890 5610
rect 7230 5550 7800 5580
rect 6150 5520 6360 5550
rect 7110 5520 7710 5550
rect 6060 5490 6360 5520
rect 7050 5490 7620 5520
rect 5970 5460 6330 5490
rect 6960 5460 7530 5490
rect 8850 5460 8910 5490
rect 5910 5430 6300 5460
rect 6870 5430 7440 5460
rect 8850 5430 8970 5460
rect 5820 5400 6210 5430
rect 6780 5400 7350 5430
rect 8880 5400 9000 5430
rect 5730 5370 6150 5400
rect 6690 5370 7290 5400
rect 8880 5370 9060 5400
rect 5610 5340 6090 5370
rect 6630 5340 7200 5370
rect 8880 5340 9120 5370
rect 5490 5310 6030 5340
rect 6540 5310 7110 5340
rect 8880 5310 9150 5340
rect 5400 5280 5940 5310
rect 6480 5280 7020 5310
rect 8880 5280 9210 5310
rect 5370 5250 5850 5280
rect 6360 5250 6960 5280
rect 8880 5250 9240 5280
rect 5340 5220 5760 5250
rect 6300 5220 6870 5250
rect 8880 5220 9270 5250
rect 9630 5220 9870 5730
rect 10110 5700 10410 5730
rect 11010 5700 11310 5730
rect 11760 5700 12210 5730
rect 10110 5670 10380 5700
rect 10080 5640 10350 5670
rect 11040 5640 11310 5700
rect 11850 5670 12240 5700
rect 11910 5640 12240 5670
rect 10080 5610 10320 5640
rect 10050 5580 10320 5610
rect 11070 5610 11310 5640
rect 10050 5520 10290 5580
rect 10020 5490 10290 5520
rect 10020 5280 10260 5490
rect 11070 5400 11340 5610
rect 11970 5460 12240 5640
rect 11580 5430 11610 5460
rect 11940 5430 12210 5460
rect 11580 5400 11640 5430
rect 11880 5400 12210 5430
rect 11070 5370 11310 5400
rect 11580 5370 12180 5400
rect 11040 5280 11310 5370
rect 11550 5340 12180 5370
rect 11550 5310 12150 5340
rect 11520 5280 12120 5310
rect 10020 5250 10290 5280
rect 11010 5250 11280 5280
rect 11490 5250 12090 5280
rect 10050 5220 10290 5250
rect 10980 5220 11280 5250
rect 11430 5220 12060 5250
rect 5340 5190 5670 5220
rect 6240 5190 6780 5220
rect 7980 5190 8280 5220
rect 8880 5190 9330 5220
rect 5370 5160 5550 5190
rect 6180 5160 6690 5190
rect 7890 5160 8370 5190
rect 8880 5160 9360 5190
rect 5400 5130 5490 5160
rect 6150 5130 6600 5160
rect 7830 5130 8430 5160
rect 8880 5130 9390 5160
rect 6120 5100 6510 5130
rect 7800 5100 8490 5130
rect 8880 5100 9420 5130
rect 6120 5070 6450 5100
rect 7740 5070 8520 5100
rect 8880 5070 9480 5100
rect 6120 5040 6360 5070
rect 7710 5040 8550 5070
rect 8880 5040 9510 5070
rect 5910 5010 6000 5040
rect 5790 4980 6000 5010
rect 5670 4950 5970 4980
rect 5580 4920 5970 4950
rect 5460 4890 5970 4920
rect 5400 4860 5940 4890
rect 5370 4830 5820 4860
rect 5340 4800 5700 4830
rect 5370 4770 5610 4800
rect 5370 4740 5520 4770
rect 5400 4710 5430 4740
rect 5880 4590 5970 4620
rect 5790 4560 5970 4590
rect 5670 4530 6000 4560
rect 5580 4500 6000 4530
rect 5460 4470 6000 4500
rect 5400 4440 5940 4470
rect 5370 4410 5820 4440
rect 5340 4380 5700 4410
rect 5370 4350 5610 4380
rect 5370 4320 5520 4350
rect 5400 4290 5430 4320
rect 5880 4170 5970 4200
rect 5790 4140 5970 4170
rect 5670 4110 5970 4140
rect 5580 4080 6000 4110
rect 5460 4050 5970 4080
rect 5400 4020 5910 4050
rect 5370 3990 5820 4020
rect 5340 3960 5730 3990
rect 5370 3930 5640 3960
rect 5370 3900 5520 3930
rect 5400 3870 5460 3900
rect 5880 3750 5970 3780
rect 5790 3720 5970 3750
rect 5670 3690 5970 3720
rect 5580 3660 6000 3690
rect 5460 3630 5970 3660
rect 5400 3600 5910 3630
rect 5370 3570 5820 3600
rect 5340 3540 5730 3570
rect 5340 3510 5640 3540
rect 5370 3480 5550 3510
rect 5400 3450 5460 3480
rect 5880 3330 5970 3360
rect 5760 3300 5970 3330
rect 5700 3270 5970 3300
rect 5580 3240 5970 3270
rect 5430 3210 5970 3240
rect 5400 3180 5880 3210
rect 5370 3150 5790 3180
rect 5340 3120 5700 3150
rect 5340 3090 5610 3120
rect 5370 3060 5520 3090
rect 6120 2880 6330 5040
rect 7680 5010 8580 5040
rect 8880 5010 9540 5040
rect 7620 4980 8610 5010
rect 7620 4950 8070 4980
rect 8190 4950 8640 4980
rect 7590 4920 7950 4950
rect 8310 4920 8640 4950
rect 7560 4890 7890 4920
rect 8370 4890 8670 4920
rect 7530 4860 7860 4890
rect 8400 4860 8670 4890
rect 7200 4830 7230 4860
rect 7530 4830 7830 4860
rect 7020 4800 7290 4830
rect 6930 4770 7290 4800
rect 7500 4770 7770 4830
rect 8430 4800 8700 4860
rect 6840 4740 7260 4770
rect 7470 4740 7740 4770
rect 6780 4710 7230 4740
rect 7470 4710 7710 4740
rect 8460 4710 8730 4800
rect 6750 4680 7230 4710
rect 7440 4680 7710 4710
rect 6690 4650 7200 4680
rect 6660 4620 7200 4650
rect 6630 4590 7200 4620
rect 6630 4560 7020 4590
rect 7050 4560 7200 4590
rect 7440 4560 7680 4680
rect 8490 4560 8730 4710
rect 6600 4530 6930 4560
rect 6570 4500 6870 4530
rect 6570 4470 6840 4500
rect 6570 4320 6810 4470
rect 7410 4440 7680 4560
rect 8460 4470 8730 4560
rect 8460 4440 8700 4470
rect 7440 4350 7680 4440
rect 8430 4380 8700 4440
rect 8400 4350 8670 4380
rect 6570 4290 6840 4320
rect 7440 4290 7710 4350
rect 8370 4320 8670 4350
rect 8340 4290 8640 4320
rect 6570 4260 6900 4290
rect 7470 4260 7740 4290
rect 8310 4260 8640 4290
rect 8880 4260 9120 5010
rect 9150 4980 9600 5010
rect 9630 4980 9900 5220
rect 10050 5160 10320 5220
rect 10980 5190 11250 5220
rect 11490 5190 12000 5220
rect 10950 5160 11250 5190
rect 11550 5160 11940 5190
rect 10080 5130 10350 5160
rect 10920 5130 11220 5160
rect 11640 5130 11880 5160
rect 10080 5100 10380 5130
rect 10860 5100 11220 5130
rect 10110 5070 10440 5100
rect 10800 5070 11190 5100
rect 12510 5070 12690 6900
rect 13380 6840 13410 6870
rect 13290 6810 13440 6840
rect 13170 6780 13470 6810
rect 13050 6750 13470 6780
rect 12930 6720 13440 6750
rect 12840 6690 13410 6720
rect 12840 6660 13320 6690
rect 12840 6630 13200 6660
rect 12840 6600 13110 6630
rect 12840 6570 12990 6600
rect 12870 6540 12900 6570
rect 13380 6450 13410 6480
rect 13290 6420 13440 6450
rect 13200 6390 13470 6420
rect 13110 6360 13470 6390
rect 12990 6330 13470 6360
rect 12870 6300 13410 6330
rect 12840 6270 13350 6300
rect 12840 6240 13230 6270
rect 12840 6210 13140 6240
rect 12870 6180 13020 6210
rect 12870 6150 12930 6180
rect 13380 6030 13410 6060
rect 13290 6000 13470 6030
rect 13200 5970 13470 6000
rect 13080 5940 13470 5970
rect 12960 5910 13470 5940
rect 12870 5880 13410 5910
rect 12840 5850 13320 5880
rect 12840 5820 13230 5850
rect 12840 5790 13110 5820
rect 12840 5760 13020 5790
rect 12870 5730 12930 5760
rect 13350 5610 13440 5640
rect 13260 5580 13470 5610
rect 13170 5550 13470 5580
rect 13050 5520 13470 5550
rect 12930 5490 13470 5520
rect 12840 5460 13410 5490
rect 12840 5430 13290 5460
rect 12840 5400 13200 5430
rect 12840 5370 13110 5400
rect 12840 5340 12990 5370
rect 12870 5310 12930 5340
rect 13320 5190 13440 5220
rect 13230 5160 13470 5190
rect 13110 5130 13470 5160
rect 13020 5100 13470 5130
rect 12870 5070 13440 5100
rect 10110 5040 10500 5070
rect 10740 5040 11160 5070
rect 10140 5010 11130 5040
rect 12480 5010 12690 5070
rect 12840 5040 13380 5070
rect 12840 5010 13260 5040
rect 10170 4980 11100 5010
rect 12450 4980 12690 5010
rect 9210 4950 9900 4980
rect 10200 4950 11070 4980
rect 12420 4950 12690 4980
rect 12870 4980 13140 5010
rect 12870 4950 13050 4980
rect 9240 4920 9900 4950
rect 10230 4920 11040 4950
rect 12300 4920 12660 4950
rect 12870 4920 12930 4950
rect 9270 4890 9900 4920
rect 10260 4890 11010 4920
rect 12210 4890 12660 4920
rect 9300 4860 9900 4890
rect 10320 4860 10950 4890
rect 12120 4860 12630 4890
rect 9360 4830 9900 4860
rect 10380 4830 10890 4860
rect 12030 4830 12600 4860
rect 9390 4800 9900 4830
rect 10440 4800 10800 4830
rect 11940 4800 12540 4830
rect 13320 4800 13410 4830
rect 9450 4770 9900 4800
rect 10590 4770 10680 4800
rect 11850 4770 12480 4800
rect 13230 4770 13440 4800
rect 9480 4740 9900 4770
rect 11760 4740 12390 4770
rect 13140 4740 13470 4770
rect 9510 4710 9900 4740
rect 11670 4710 12330 4740
rect 13050 4710 13470 4740
rect 9570 4680 9900 4710
rect 11580 4680 12240 4710
rect 12930 4680 13440 4710
rect 9600 4650 9900 4680
rect 11490 4650 12120 4680
rect 12720 4650 12780 4680
rect 12870 4650 13380 4680
rect 9630 4620 9900 4650
rect 11400 4620 12030 4650
rect 12630 4620 12750 4650
rect 9690 4590 9900 4620
rect 11310 4590 11970 4620
rect 12600 4590 12750 4620
rect 9720 4560 9900 4590
rect 11250 4560 11850 4590
rect 12570 4560 12750 4590
rect 12870 4620 13290 4650
rect 12870 4590 13200 4620
rect 12870 4560 13110 4590
rect 9780 4530 9900 4560
rect 11160 4530 11760 4560
rect 12570 4530 12720 4560
rect 9810 4500 9900 4530
rect 11040 4500 11670 4530
rect 10980 4470 11580 4500
rect 12240 4470 12270 4500
rect 12540 4470 12720 4530
rect 12870 4530 12990 4560
rect 12870 4500 12930 4530
rect 10890 4440 11520 4470
rect 12180 4440 12300 4470
rect 10800 4410 11430 4440
rect 12060 4410 12300 4440
rect 10710 4380 11340 4410
rect 11970 4380 12300 4410
rect 12510 4410 12690 4470
rect 12510 4380 12660 4410
rect 10620 4350 11250 4380
rect 11910 4350 12060 4380
rect 12090 4350 12330 4380
rect 10530 4320 11160 4350
rect 11820 4320 12060 4350
rect 12120 4320 12360 4350
rect 10440 4290 11070 4320
rect 11730 4290 12090 4320
rect 10380 4260 10980 4290
rect 11640 4260 12090 4290
rect 12150 4290 12360 4320
rect 12480 4320 12660 4380
rect 12480 4290 12630 4320
rect 12150 4260 12390 4290
rect 6600 4230 6960 4260
rect 7470 4230 7770 4260
rect 8280 4230 8610 4260
rect 8880 4230 9090 4260
rect 10290 4230 10890 4260
rect 11550 4230 12060 4260
rect 12180 4230 12390 4260
rect 12450 4260 12630 4290
rect 12450 4230 12600 4260
rect 6600 4200 7050 4230
rect 7500 4200 7800 4230
rect 8220 4200 8580 4230
rect 8910 4200 8970 4230
rect 10200 4200 10800 4230
rect 11520 4200 12000 4230
rect 12210 4200 12600 4230
rect 6630 4170 7170 4200
rect 7500 4170 7860 4200
rect 8160 4170 8550 4200
rect 10110 4170 10710 4200
rect 6660 4140 7230 4170
rect 7530 4140 7950 4170
rect 8070 4140 8550 4170
rect 10020 4140 10650 4170
rect 6690 4110 7290 4140
rect 7560 4110 8520 4140
rect 9930 4110 10560 4140
rect 11520 4110 11910 4200
rect 12210 4170 12570 4200
rect 12240 4140 12570 4170
rect 6720 4080 7320 4110
rect 7590 4080 8490 4110
rect 9870 4080 10470 4110
rect 11160 4080 11280 4110
rect 11520 4080 11670 4110
rect 6780 4050 7350 4080
rect 7620 4050 8460 4080
rect 9780 4050 10380 4080
rect 11070 4050 11340 4080
rect 11520 4050 11580 4080
rect 6840 4020 7350 4050
rect 7650 4020 8400 4050
rect 9690 4020 10290 4050
rect 10980 4020 11400 4050
rect 6930 3990 7350 4020
rect 7710 3990 8370 4020
rect 9600 3990 10200 4020
rect 10920 3990 11430 4020
rect 7020 3960 7380 3990
rect 7770 3960 8310 3990
rect 9510 3960 10140 3990
rect 7110 3870 7380 3960
rect 7830 3930 8250 3960
rect 9420 3930 10050 3960
rect 10890 3930 11460 3990
rect 7920 3900 8160 3930
rect 9330 3900 9960 3930
rect 10890 3900 11490 3930
rect 9240 3870 9870 3900
rect 10890 3870 11100 3900
rect 7110 3840 7350 3870
rect 9150 3840 9780 3870
rect 7080 3780 7350 3840
rect 9090 3810 9690 3840
rect 9000 3780 9600 3810
rect 7050 3750 7320 3780
rect 8910 3750 9510 3780
rect 10410 3750 10470 3810
rect 6690 3720 6780 3750
rect 6990 3720 7320 3750
rect 8820 3720 9420 3750
rect 10380 3720 10500 3750
rect 6690 3690 7290 3720
rect 8730 3690 9330 3720
rect 10380 3690 10530 3720
rect 6660 3660 7260 3690
rect 8640 3660 9240 3690
rect 10380 3660 10560 3690
rect 6630 3630 7230 3660
rect 8550 3630 9150 3660
rect 10350 3630 10560 3660
rect 10890 3630 11070 3870
rect 11280 3840 11490 3900
rect 11310 3780 11490 3840
rect 11280 3690 11460 3780
rect 11250 3660 11430 3690
rect 11190 3630 11400 3660
rect 6630 3600 7200 3630
rect 8460 3600 9090 3630
rect 9780 3600 9930 3630
rect 6600 3570 7140 3600
rect 8370 3570 9000 3600
rect 9690 3570 10020 3600
rect 10350 3570 10590 3630
rect 10890 3600 11400 3630
rect 10890 3570 11370 3600
rect 6570 3540 7110 3570
rect 8280 3540 8910 3570
rect 9600 3540 10050 3570
rect 6570 3510 7050 3540
rect 8190 3510 8820 3540
rect 9540 3510 10080 3540
rect 10320 3510 10620 3570
rect 10890 3540 11340 3570
rect 10890 3510 11310 3540
rect 6660 3480 6990 3510
rect 8100 3480 8760 3510
rect 8010 3450 8640 3480
rect 9510 3450 10110 3510
rect 10290 3480 10650 3510
rect 10890 3480 11340 3510
rect 11730 3480 11910 4110
rect 12270 4080 12540 4140
rect 12300 4050 12540 4080
rect 12330 4020 12540 4050
rect 12330 3810 12510 4020
rect 12330 3750 12540 3810
rect 12330 3720 12510 3750
rect 12360 3690 12480 3720
rect 12360 3660 12390 3690
rect 10290 3450 10680 3480
rect 7920 3420 8550 3450
rect 9510 3420 9810 3450
rect 9870 3420 10140 3450
rect 7860 3390 8460 3420
rect 7770 3360 8400 3390
rect 9090 3360 9150 3390
rect 7680 3330 8310 3360
rect 9000 3330 9150 3360
rect 7590 3300 8190 3330
rect 7500 3270 8130 3300
rect 7410 3240 8040 3270
rect 7320 3210 7920 3240
rect 7230 3180 7860 3210
rect 8610 3180 8700 3210
rect 7140 3150 7770 3180
rect 8550 3150 8700 3180
rect 7050 3120 7680 3150
rect 6960 3090 7620 3120
rect 6870 3060 7530 3090
rect 8520 3060 8700 3150
rect 6780 3030 7410 3060
rect 6690 3000 7320 3030
rect 8100 3000 8310 3030
rect 6600 2970 7230 3000
rect 8040 2970 8370 3000
rect 6540 2940 7170 2970
rect 8010 2940 8400 2970
rect 6450 2910 7080 2940
rect 7980 2910 8400 2940
rect 6360 2880 6990 2910
rect 7950 2880 8370 2910
rect 6120 2850 6870 2880
rect 7950 2850 8340 2880
rect 8550 2850 8700 3060
rect 8970 3150 9150 3330
rect 9510 3240 9720 3420
rect 9930 3300 10140 3420
rect 10260 3390 10680 3450
rect 10890 3450 11400 3480
rect 11730 3450 11880 3480
rect 10890 3420 11100 3450
rect 11160 3420 11430 3450
rect 11760 3420 11790 3450
rect 10260 3360 10440 3390
rect 10230 3330 10440 3360
rect 10500 3330 10710 3390
rect 10230 3300 10410 3330
rect 10530 3300 10740 3330
rect 9930 3240 10110 3300
rect 9510 3150 9690 3240
rect 9900 3210 10110 3240
rect 10200 3270 10410 3300
rect 10200 3210 10380 3270
rect 10560 3240 10770 3300
rect 10470 3210 10800 3240
rect 9870 3180 10080 3210
rect 10170 3180 10800 3210
rect 10890 3180 11070 3420
rect 11190 3390 11460 3420
rect 11220 3360 11490 3390
rect 11250 3330 11520 3360
rect 11280 3300 11490 3330
rect 12000 3300 12120 3330
rect 11310 3270 11400 3300
rect 11970 3270 12150 3300
rect 9780 3150 10050 3180
rect 10170 3150 10830 3180
rect 8970 2940 9180 3150
rect 8910 2910 9180 2940
rect 8820 2880 9180 2910
rect 8730 2850 9180 2880
rect 6120 2820 6810 2850
rect 7920 2820 8130 2850
rect 8220 2820 8310 2850
rect 6120 2790 6690 2820
rect 6120 2760 6600 2790
rect 6120 2730 6540 2760
rect 7470 2730 7500 2790
rect 6120 2700 6450 2730
rect 7440 2700 7530 2730
rect 7890 2700 8070 2820
rect 8550 2760 9180 2850
rect 8550 2730 8910 2760
rect 9000 2730 9180 2760
rect 8550 2700 8820 2730
rect 6120 2670 6360 2700
rect 6120 2640 6300 2670
rect 7440 2640 7560 2700
rect 7890 2670 8100 2700
rect 7890 2640 8220 2670
rect 6120 2610 6210 2640
rect 7410 2580 7590 2640
rect 7890 2610 8340 2640
rect 7920 2580 8370 2610
rect 6780 2550 6810 2580
rect 6690 2520 6810 2550
rect 6660 2460 6810 2520
rect 7380 2550 7620 2580
rect 7950 2550 8400 2580
rect 8550 2550 8730 2700
rect 7380 2490 7650 2550
rect 7980 2520 8430 2550
rect 8040 2490 8430 2520
rect 6450 2430 6570 2460
rect 6360 2400 6570 2430
rect 6270 2370 6570 2400
rect 6210 2340 6570 2370
rect 6120 2310 6570 2340
rect 6090 2280 6570 2310
rect 6090 2250 6540 2280
rect 6090 2220 6420 2250
rect 6090 2190 6330 2220
rect 6090 2010 6270 2190
rect 6420 2040 6510 2070
rect 6330 2010 6510 2040
rect 6090 1920 6540 2010
rect 6090 1890 6510 1920
rect 6090 1860 6450 1890
rect 6660 1860 6840 2460
rect 7350 2430 7680 2490
rect 8190 2460 8460 2490
rect 7350 2400 7710 2430
rect 7320 2370 7740 2400
rect 7320 2310 7500 2370
rect 7530 2340 7740 2370
rect 8250 2370 8460 2460
rect 8250 2340 8430 2370
rect 7320 2280 7470 2310
rect 7560 2280 7770 2340
rect 8010 2310 8040 2340
rect 8220 2310 8430 2340
rect 8520 2310 8730 2550
rect 8970 2490 9180 2730
rect 9510 3120 10020 3150
rect 10140 3120 10830 3150
rect 10890 3150 11040 3180
rect 10890 3120 10950 3150
rect 9510 3090 9990 3120
rect 10140 3090 10560 3120
rect 10620 3090 10830 3120
rect 9510 3060 9960 3090
rect 10110 3060 10470 3090
rect 10650 3060 10770 3090
rect 9510 3030 9930 3060
rect 10110 3030 10380 3060
rect 10650 3030 10680 3060
rect 12000 3030 12150 3270
rect 9510 3000 9870 3030
rect 9510 2970 9780 3000
rect 10080 2970 10290 3030
rect 9510 2700 9690 2970
rect 10050 2880 10260 2970
rect 10020 2850 10200 2880
rect 10020 2820 10080 2850
rect 12000 2760 12180 3030
rect 11880 2730 12300 2760
rect 11820 2700 12360 2730
rect 9510 2670 9660 2700
rect 11760 2670 12420 2700
rect 9540 2640 9570 2670
rect 11730 2640 12450 2670
rect 11700 2610 12480 2640
rect 11670 2580 11970 2610
rect 12210 2580 12510 2610
rect 11640 2550 11910 2580
rect 12300 2550 12540 2580
rect 11640 2520 11850 2550
rect 12360 2520 12570 2550
rect 11610 2490 11820 2520
rect 12390 2490 12600 2520
rect 9000 2460 9150 2490
rect 9000 2430 9030 2460
rect 11580 2430 11790 2490
rect 12420 2460 12600 2490
rect 12420 2430 12630 2460
rect 11550 2400 11760 2430
rect 12000 2400 12210 2430
rect 12450 2400 12630 2430
rect 11550 2370 11730 2400
rect 11970 2370 12240 2400
rect 11520 2340 11730 2370
rect 11940 2340 12300 2370
rect 7980 2280 8400 2310
rect 8520 2280 8670 2310
rect 7290 2220 7470 2280
rect 7590 2220 7800 2280
rect 7950 2250 8400 2280
rect 8550 2250 8580 2280
rect 11520 2250 11700 2340
rect 11910 2310 12300 2340
rect 12480 2310 12660 2400
rect 11880 2280 12060 2310
rect 12150 2280 12330 2310
rect 7920 2220 8370 2250
rect 7290 2190 7440 2220
rect 7590 2190 7830 2220
rect 7890 2190 8340 2220
rect 7260 2160 7440 2190
rect 7530 2160 7860 2190
rect 7920 2160 8310 2190
rect 7260 2100 7890 2160
rect 7950 2130 8280 2160
rect 8010 2100 8220 2130
rect 11490 2100 11700 2250
rect 11850 2250 12030 2280
rect 12180 2250 12330 2280
rect 11850 2130 12000 2250
rect 12210 2130 12360 2250
rect 11850 2100 12030 2130
rect 12180 2100 12330 2130
rect 7230 2070 7920 2100
rect 7230 2040 7620 2070
rect 7710 2040 7950 2070
rect 7230 2010 7560 2040
rect 7710 2010 7920 2040
rect 11520 2010 11700 2100
rect 11880 2070 12330 2100
rect 12510 2070 12690 2310
rect 11880 2040 12300 2070
rect 12480 2040 12690 2070
rect 11910 2010 12270 2040
rect 7200 1980 7470 2010
rect 7740 1980 7800 2010
rect 11520 1980 11730 2010
rect 11940 1980 12240 2010
rect 12480 1980 12660 2040
rect 7200 1950 7380 1980
rect 11550 1950 11730 1980
rect 12000 1950 12210 1980
rect 12450 1950 12660 1980
rect 7170 1920 7350 1950
rect 11550 1920 11760 1950
rect 7020 1890 7350 1920
rect 6900 1860 7350 1890
rect 11580 1890 11790 1920
rect 12420 1890 12630 1950
rect 11580 1860 11820 1890
rect 12390 1860 12600 1890
rect 6090 1830 6360 1860
rect 6660 1830 7350 1860
rect 11610 1830 11850 1860
rect 12330 1830 12570 1860
rect 6090 1800 6300 1830
rect 6660 1800 7320 1830
rect 11640 1800 11910 1830
rect 12270 1800 12540 1830
rect 6090 1410 6270 1800
rect 6660 1770 7200 1800
rect 11670 1770 12000 1800
rect 12210 1770 12510 1800
rect 6660 1740 7110 1770
rect 11700 1740 12480 1770
rect 6660 1710 7050 1740
rect 11730 1710 12450 1740
rect 6660 1680 6960 1710
rect 11760 1680 12420 1710
rect 6660 1650 6870 1680
rect 11820 1650 12360 1680
rect 6660 1620 6780 1650
rect 11880 1620 12300 1650
rect 6660 1590 6690 1620
rect 11970 1590 12210 1620
rect 6090 1380 6180 1410
<< end >>
