magic
tech sky130A
magscale 1 2
timestamp 1740521415
<< error_s >>
rect 9308 28387 9352 28477
<< metal2 >>
rect 4716 36006 5116 36016
rect 4716 35596 5116 35606
rect 4852 33660 5068 33670
rect 4852 33454 5068 33464
rect 4810 29448 5186 29458
rect 4810 29038 5186 29048
rect 13944 28352 14012 28362
rect 13944 28274 14012 28284
rect 4776 27872 5128 27882
rect 4776 27486 5128 27496
rect 4868 27152 5012 27162
rect 4868 26996 5012 27006
rect 18756 26014 18916 26024
rect 18756 25894 18916 25904
rect 18206 25836 18316 25846
rect 18206 25712 18316 25722
rect 7386 25250 7566 25260
rect 7386 25060 7566 25070
<< via2 >>
rect 4716 35606 5116 36006
rect 4852 33464 5068 33660
rect 4810 29048 5186 29448
rect 13944 28284 14012 28352
rect 4776 27496 5128 27872
rect 4868 27006 5012 27152
rect 18756 25904 18916 26014
rect 18206 25722 18316 25836
rect 7386 25070 7566 25250
<< metal3 >>
rect 4706 36006 5126 36011
rect 4706 35606 4716 36006
rect 5116 35606 5126 36006
rect 4706 35601 5126 35606
rect 4842 33660 5078 33665
rect 4842 33464 4852 33660
rect 5068 33464 5078 33660
rect 4842 33459 5078 33464
rect 804 29040 814 29464
rect 1164 29448 5210 29464
rect 1164 29048 4810 29448
rect 5186 29048 5210 29448
rect 1164 29040 5210 29048
rect 13906 28352 14036 28410
rect 13906 28284 13944 28352
rect 14012 28284 14036 28352
rect 13906 28254 14036 28284
rect 206 27488 216 27896
rect 568 27888 578 27896
rect 568 27872 5152 27888
rect 568 27496 4776 27872
rect 5128 27496 5152 27872
rect 568 27488 5152 27496
rect 4858 27152 5022 27157
rect 4858 27006 4868 27152
rect 5012 27006 5022 27152
rect 4858 27001 5022 27006
rect 18746 26014 18926 26019
rect 18746 25904 18756 26014
rect 18916 25904 18926 26014
rect 18746 25899 18926 25904
rect 18196 25836 18326 25841
rect 18196 25722 18206 25836
rect 18316 25722 18326 25836
rect 18196 25717 18326 25722
rect 7376 25250 7576 25255
rect 7376 25070 7386 25250
rect 7566 25070 7576 25250
rect 7376 25065 7576 25070
<< via3 >>
rect 4716 35606 5116 36006
rect 4852 33464 5068 33660
rect 814 29040 1164 29464
rect 13944 28284 14012 28352
rect 216 27488 568 27896
rect 4868 27006 5012 27152
rect 18756 25904 18916 26014
rect 18206 25722 18316 25836
rect 7386 25070 7566 25250
<< metal4 >>
rect 3006 44990 3066 45152
rect 3558 44990 3618 45152
rect 4110 44990 4170 45152
rect 4662 44990 4722 45152
rect 5214 44990 5274 45152
rect 5766 44990 5826 45152
rect 6318 44990 6378 45152
rect 6870 44990 6930 45152
rect 7422 44990 7482 45152
rect 7974 44990 8034 45152
rect 8526 44990 8586 45152
rect 9078 44990 9138 45152
rect 9630 44990 9690 45152
rect 10182 44990 10242 45152
rect 10734 44990 10794 45152
rect 11286 44990 11346 45152
rect 11838 44990 11898 45152
rect 12390 44990 12450 45152
rect 12942 44990 13002 45152
rect 13494 44990 13554 45152
rect 14046 44990 14106 45152
rect 14598 44990 14658 45152
rect 15150 44990 15210 45152
rect 922 44842 15212 44990
rect 922 44152 1070 44842
rect 200 27896 600 44152
rect 200 27488 216 27896
rect 568 27488 600 27896
rect 200 1000 600 27488
rect 800 29464 1200 44152
rect 800 29040 814 29464
rect 1164 29040 1200 29464
rect 800 1000 1200 29040
rect 1400 36006 1800 44152
rect 15702 42078 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 15702 42018 23046 42078
rect 4715 36006 5117 36007
rect 1400 35606 4716 36006
rect 5116 35606 5117 36006
rect 1400 1000 1800 35606
rect 4715 35605 5117 35606
rect 4851 33660 5069 33661
rect 4851 33570 4852 33660
rect 4686 33510 4852 33570
rect 4686 25650 4746 33510
rect 4851 33464 4852 33510
rect 5068 33464 5069 33660
rect 4851 33463 5069 33464
rect 22986 29482 23046 42018
rect 13948 29422 23046 29482
rect 13948 28353 14008 29422
rect 13943 28352 14013 28353
rect 13943 28284 13944 28352
rect 14012 28284 14013 28352
rect 13943 28283 14013 28284
rect 4867 27152 5013 27153
rect 4867 27006 4868 27152
rect 5012 27006 5013 27152
rect 4867 27005 5013 27006
rect 4910 26308 4970 27005
rect 23430 26308 23490 45152
rect 4910 26248 23490 26308
rect 18755 26014 18917 26015
rect 18755 25904 18756 26014
rect 18916 25992 18917 26014
rect 23982 25992 24042 45152
rect 18916 25932 24042 25992
rect 18916 25904 18917 25932
rect 18755 25903 18917 25904
rect 18205 25836 18317 25837
rect 18205 25722 18206 25836
rect 18316 25812 18317 25836
rect 24534 25812 24594 45152
rect 25086 44952 25146 45152
rect 18316 25752 24594 25812
rect 18316 25722 18317 25752
rect 18205 25721 18317 25722
rect 25638 25650 25698 45152
rect 26190 44952 26250 45152
rect 4686 25590 25698 25650
rect 7385 25250 7567 25251
rect 7385 25070 7386 25250
rect 7566 25070 7567 25250
rect 7385 25069 7567 25070
rect 7386 23478 7566 25069
rect 7386 23298 27414 23478
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 0 27414 23298
use flash  flash_0 flash
timestamp 1740521415
transform 1 0 4812 0 1 25950
box -103 -1220 18127 15751
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 1400 1000 1800 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
