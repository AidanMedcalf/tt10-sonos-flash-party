** sch_path: /home/uri/p/tt10-sonos-flash-party/xschem/level_shifter_tb.sch
**.subckt level_shifter_tb
V1 VPROG GND 10
V2 clk GND PULSE(0 1.8 0 0 0 250n 500n)
V3 VDPWR GND 1.8
x4 VPROG VDPWR clk vout net1 GND GND level_shifter
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/uri/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt





.tran 10n 1u
.save all

.control
run
write level_shifter_tb.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  level_shifter.sym # of pins=7
** sym_path: /home/uri/p/tt10-sonos-flash-party/xschem/level_shifter.sym
** sch_path: /home/uri/p/tt10-sonos-flash-party/xschem/level_shifter.sch
.subckt level_shifter avdd dvdd in out out_b avss dvss
*.iopin avdd
*.opin out_b
*.opin out
*.iopin avss
*.iopin dvdd
*.ipin in
*.iopin dvss
XM1 in_b in dvss dvss sky130_fd_pr__nfet_01v8 L=3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 in_b in dvdd dvdd sky130_fd_pr__pfet_01v8 L=3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 out_b out avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 out out_b avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 out in_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=3 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 out_b in avss avss sky130_fd_pr__nfet_g5v0d10v5 L=3 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XD3 dvss in sky130_fd_pr__diode_pw2nd_05v5 area=0.315e12 perim=4e6
.ends

.GLOBAL GND
.GLOBAL VPROG
.GLOBAL VDPWR
.end
