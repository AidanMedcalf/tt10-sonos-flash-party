* NGSPICE file created from charge_pump.ext - technology: sky130A

.subckt charge_pump VAPWR VOUT clk VGND
X0 clkina clkinb VAPWR.t4 VAPWR.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X1 clkinb clk.t0 VGND.t2 VGND.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X2 stage1 VAPWR.t7 VAPWR.t9 VAPWR.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 stage2 stage1 stage1 stage1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 clkb clkinb VGND.t8 VGND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X5 clkb clkinb VAPWR.t2 VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X6 VOUT VGND.t0 sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X7 VOUT.t0 stage2 stage2 stage2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X8 clkinb clk.t1 VAPWR.t6 VAPWR.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X9 clkina clkinb VGND.t6 VGND.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X10 clka clkina VGND.t4 VGND.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X11 clka clkina VAPWR.t1 VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X12 clkb stage2 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X13 clka stage1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
R0 VAPWR.n0 VAPWR.t3 28.5727
R1 VAPWR.t5 VAPWR 355.541
R2 VAPWR.n5 VAPWR.n2 1577.4
R3 VAPWR.n8 VAPWR.n4 1577.4
R4 VAPWR.n6 VAPWR.n4 722.497
R5 VAPWR.n7 VAPWR.n2 722.497
R6 VAPWR VAPWR.t4 649.99
R7 VAPWR VAPWR.t6 649.765
R8 VAPWR.t5 VAPWR.t3 487.901
R9 VAPWR VAPWR.t7 236.188
R10 VAPWR.t7 VAPWR 236.011
R11 VAPWR VAPWR.n3 184.847
R12 VAPWR.n3 VAPWR.n1 184.847
R13 VAPWR VAPWR.t2 167.41
R14 VAPWR VAPWR.t1 167.19
R15 VAPWR VAPWR.n8 146.25
R16 VAPWR.n5 VAPWR.n1 146.25
R17 VAPWR VAPWR.n2 98.9887
R18 VAPWR.n4 VAPWR.n3 97.5005
R19 VAPWR.n0 VAPWR.t0 3.34151
R20 VAPWR VAPWR.t9 78.1972
R21 VAPWR.n6 VAPWR.n5 72.5386
R22 VAPWR.n8 VAPWR.n7 72.5386
R23 VAPWR.n7 VAPWR.t8 66.988
R24 VAPWR.t8 VAPWR.n6 66.988
R25 VAPWR VAPWR.n0 38.6117
R26 VAPWR VAPWR.n9 33.1299
R27 VAPWR VAPWR.n1 11.7843
R28 clk clk.t1 54.3383
R29 clk clk.t0 53.1307
R30 VGND.n10 VGND.n8 17010.2
R31 VGND.n3 VGND.n8 17010.2
R32 VGND.n14 VGND.n12 9438.3
R33 VGND.n20 VGND.n12 5607.68
R34 VGND.n12 VGND.n11 4686.84
R35 VGND.n18 VGND.n0 3790.36
R36 VGND.n15 VGND.n0 3790.36
R37 VGND.n11 VGND.n9 3370.76
R38 VGND.n21 VGND.n20 2547.06
R39 VGND.n21 VGND.n9 2166.87
R40 VGND.n9 VGND.n8 1472.95
R41 VGND.n4 VGND.n5 7.29093
R42 VGND.n20 VGND.n19 957.745
R43 VGND.t3 VGND.t7 838.864
R44 VGND.t1 VGND.t5 838.864
R45 VGND.n19 VGND.t7 530.34
R46 VGND.n14 VGND.t1 530.34
R47 VGND.n2 VGND.n1 0.871201
R48 VGND.n13 VGND.t3 419.433
R49 VGND.t5 VGND.n13 419.433
R50 VGND.n1 VGND.n17 267.295
R51 VGND.n1 VGND.t6 227.643
R52 VGND.n7 VGND.t2 227.398
R53 VGND.n17 VGND.n16 170.542
R54 VGND.n19 VGND.n18 97.5005
R55 VGND.n16 VGND.n15 97.5005
R56 VGND.n15 VGND.n14 97.5005
R57 VGND.n1 VGND.t4 82.9558
R58 VGND.n8 VGND.n5 27.0289
R59 VGND.n1 VGND.n0 24.3755
R60 VGND.n13 VGND.n0 24.3755
R61 VGND.n4 VGND.n3 9.28621
R62 VGND.n3 VGND.n21 9.28621
R63 VGND.n10 VGND.n6 9.28621
R64 VGND.n11 VGND.n10 9.28621
R65 VGND.n6 VGND.n5 8.15439
R66 VGND.n6 VGND 5.97887
R67 VGND.n4 VGND 5.15194
R68 VGND.n4 VGND.t0 4.15891
R69 VGND.n7 VGND.n4 4.09497
R70 VGND.n18 VGND.n2 100.788
R71 VGND.n16 VGND.n7 1.5505
R72 VGND.n7 VGND.n1 1.01429
R73 VGND.n2 VGND.t8 83.1878
R74 VOUT VOUT.t0 78.1972
R75 VOUT VOUT.n0 33.1299
C0 clkb stage2 59.0307f
C1 stage2 stage1 5.8896f
C2 clka stage1 57.614f
C3 VAPWR stage1 2.72272f
C4 VOUT VGND 72.02551f
C5 VAPWR VGND 16.19416f
C6 clkb VGND 4.70804f
C7 clka VGND 5.28435f
C8 clkinb VGND 3.10612f
C9 stage2 VGND 24.3838f
C10 stage1 VGND 22.4378f
.ends

