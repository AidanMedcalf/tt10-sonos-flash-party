* NGSPICE file created from tt_um_sonos_flash_party.ext - technology: sky130A

.subckt tt_um_sonos_flash_party clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VDPWR VGND VAPWR
X0 flash_0.x7.VPRGNEG VGND.t42 sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X1 flash_0.x7.VPRGPOS.t29 flash_0.x7.pos_mid_b.t5 flash_0.x7.vintp flash_0.x7.VPRGPOS.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X2 flash_0.x2.clkb.t0 flash_0.x2.clkinb VAPWR.t8 VAPWR.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X3 flash_0.x7.VPRGPOS.t30 flash_0.x7.pos_mid flash_0.x7.pos_mid_b.t3 flash_0.x7.VPRGPOS.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X4 flash_0.x3.clkinb clk.t0 VAPWR.t16 VAPWR.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X5 flash_0.x7.VPRGPOS.t3 flash_0.x4.pos_mid flash_0.x4.pos_mid_b.t0 flash_0.x7.VPRGPOS.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X6 VGND.t5 ui_in[1].t0 flash_0.x4.neg_en_b.t3 VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X7 flash_0.x4.dcgint.t11 flash_0.x4.neg_mid_b.t7 flash_0.x4.VOUT flash_0.x4.dcgint.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X8 flash_0.x7.pos_mid_b.t0 ui_in[1].t1 VGND.t13 VGND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X9 flash_0.x7.pos_mid flash_0.x7.pos_en_b.t4 VGND.t8 VGND.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X10 VDPWR.t43 ui_in[1].t2 flash_0.x4.neg_mid VDPWR.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X11 ua[0].t3 VGND.t40 VGND.t41 ua[0].t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=10
X12 VDPWR.t4 flash_0.x7.neg_en_b.t4 flash_0.x7.neg_mid_b.t5 VDPWR.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X13 VDPWR.t21 flash_0.x7.neg_en_b.t5 flash_0.x7.neg_mid_b.t4 VDPWR.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X14 flash_0.x5.A.t3 flash_0.x6.Y VDPWR.t52 VDPWR.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
X15 flash_0.x7.vintp flash_0.x7.pos_mid_b.t6 flash_0.x7.VPRGPOS.t28 flash_0.x7.VPRGPOS.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X16 flash_0.x7.neg_mid ui_in[0].t0 VDPWR.t18 VDPWR.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X17 flash_0.x4.neg_mid_b.t0 flash_0.x4.neg_mid flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=1
X18 flash_0.x2.clkina flash_0.x2.clkinb VAPWR.t6 VAPWR.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X19 flash_0.x4.neg_mid_b.t5 flash_0.x4.neg_en_b.t4 VDPWR.t50 VDPWR.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X20 flash_0.x7.pos_mid_b.t2 ui_in[1].t3 VGND.t36 VGND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X21 flash_0.x7.pos_mid flash_0.x7.pos_en_b.t4 VGND.t7 VGND.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X22 flash_0.x4.dcgint.t10 flash_0.x4.neg_mid_b.t8 flash_0.x4.VOUT flash_0.x4.dcgint.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X23 a_9352_28387# flash_0.x4.VOUT a_7463_28281# flash_0.x7.VOUT.t0 sky130_fd_bs_flash__special_sonosfet_star ad=0.13725 pd=1.51 as=0.13725 ps=1.51 w=0.45 l=0.22
X24 VGND.t15 ui_in[1].t4 flash_0.x7.pos_mid_b.t1 VGND.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X25 VGND.t11 ui_in[0].t1 flash_0.x4.pos_mid_b VGND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X26 flash_0.x7.VPRGNEG flash_0.x4.neg_mid_b.t9 flash_0.x4.neg_mid flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.145 ps=1.58 w=0.5 l=1
X27 flash_0.x4.vintp flash_0.x4.VDPWR1 flash_0.x4.VOUT flash_0.x7.VPRGPOS.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X28 VDPWR.t41 ui_in[1].t5 flash_0.x4.neg_en_b.t0 VDPWR.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X29 flash_0.x4.VOUT VDPWR.t58 a_16296_28578# flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X30 VDPWR.t2 flash_0.x7.neg_en_b.t6 flash_0.x7.neg_mid_b.t3 VDPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X31 w_7728_24730.t1 ua[0].t0 ua[0].t1 w_7728_24730.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
X32 flash_0.x3.stage1 VAPWR.t2 VAPWR.t4 VAPWR.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X33 flash_0.x4.VOUT flash_0.x4.VDPWR1 flash_0.x4.vintp flash_0.x7.VPRGPOS.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X34 flash_0.x7.neg_en_b.t2 ui_in[0].t2 VGND.t39 VGND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X35 flash_0.x7.pos_en_b.t3 ui_in[1].t6 VGND.t19 VGND.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X36 VGND.t70 ui_in[1].t7 flash_0.x7.pos_mid_b.t4 VGND.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X37 flash_0.x3.clka.t0 flash_0.x3.clkina VAPWR.t14 VAPWR.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X38 VGND.t10 ui_in[0].t3 flash_0.x4.pos_mid_b VGND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X39 flash_0.x3.clkb.t1 flash_0.x3.clkinb VGND.t50 VGND.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X40 flash_0.x4.vintp flash_0.x4.pos_mid_b.t3 flash_0.x7.VPRGPOS.t32 flash_0.x7.VPRGPOS.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X41 flash_0.x4.VOUT VDPWR.t59 a_16296_28578# flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X42 flash_0.x4.dcgint.t2 flash_0.x4.pos_en_b.t4 VGND.t58 VGND.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X43 flash_0.x7.VPRGPOS.t5 flash_0.x4.pos_mid_b.t4 flash_0.x4.vintp flash_0.x7.VPRGPOS.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X44 flash_0.x6.Y ui_in[2].t0 VGND.t63 VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X45 flash_0.x7.VOUT.t6 flash_0.x7.VDPWR1 flash_0.x7.vintp flash_0.x7.VPRGPOS.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X46 flash_0.x2.clka.t1 flash_0.x2.clkina VGND.t52 VGND.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X47 flash_0.x3.clkb flash_0.x3.stage2 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X48 VGND.t24 ui_in[1].t8 flash_0.x7.pos_en_b.t2 VGND.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X49 VGND.t38 ui_in[0].t4 flash_0.x4.pos_en_b.t3 VGND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X50 VDPWR.t49 flash_0.x4.neg_en_b.t5 flash_0.x4.neg_mid_b.t4 VDPWR.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X51 flash_0.x7.neg_en_b.t0 ui_in[0].t5 VDPWR.t8 VDPWR.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=3
X52 flash_0.x7.pos_en_b.t0 ui_in[1].t9 VDPWR.t39 VDPWR.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X53 flash_0.x4.dcgint.t1 flash_0.x4.pos_en_b.t4 VGND.t56 VGND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X54 VDPWR.t37 ui_in[1].t10 flash_0.x4.neg_mid VDPWR.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X55 a_16296_28578# flash_0.x4.neg_mid_b.t10 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X56 flash_0.x4.neg_mid_b.t2 flash_0.x4.neg_en_b.t6 VDPWR.t48 VDPWR.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X57 flash_0.x7.VPRGPOS.t27 flash_0.x7.pos_mid_b.t7 flash_0.x7.vintp flash_0.x7.VPRGPOS.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X58 flash_0.x7.neg_mid ui_in[0].t6 VDPWR.t57 VDPWR.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X59 flash_0.x4.neg_mid_b.t6 flash_0.x4.neg_en_b.t7 VDPWR.t47 VDPWR.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X60 flash_0.x4.dcgint.t8 flash_0.x4.neg_mid_b.t11 flash_0.x4.VOUT flash_0.x4.dcgint.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X61 flash_0.x7.VPRGPOS.t1 w_7728_24730.t2 w_7728_24730.t3 flash_0.x7.VPRGPOS.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
X62 VDPWR.t35 ui_in[1].t11 flash_0.x7.pos_en_b.t1 VDPWR.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X63 flash_0.x3.clkinb clk.t1 VGND.t21 VGND.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X64 VDPWR.t56 ui_in[0].t7 flash_0.x4.pos_en_b.t1 VDPWR.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X65 flash_0.x2.clkina flash_0.x2.clkinb VGND.t46 VGND.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X66 flash_0.x3.clka flash_0.x3.stage1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X67 a_16296_28578# flash_0.x4.neg_mid_b.t10 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X68 flash_0.x4.dcgint.t0 flash_0.x4.pos_en_b.t4 VGND.t54 VGND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X69 flash_0.x4.VOUT flash_0.x4.neg_mid_b.t12 flash_0.x4.dcgint.t7 flash_0.x4.dcgint.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X70 flash_0.x4.dcgint.t6 flash_0.x4.neg_mid_b.t13 flash_0.x4.VOUT flash_0.x4.dcgint.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X71 flash_0.x4.vintp flash_0.x4.VDPWR1 flash_0.x4.VOUT flash_0.x7.VPRGPOS.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X72 a_7463_28281# ui_in[2].t1 VGND.t60 VGND.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X73 flash_0.x7.neg_mid ui_in[0].t8 VDPWR.t17 VDPWR.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X74 flash_0.x7.dcgint.t8 flash_0.x7.neg_mid_b.t7 flash_0.x7.VOUT.t11 flash_0.x7.dcgint.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X75 VDPWR.t44 ui_in[0].t9 flash_0.x7.neg_mid VDPWR.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X76 uo_out[0].t0 flash_0.x5.A.t4 VDPWR.t20 VDPWR.t19 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X77 VDPWR.t6 ui_in[0].t10 flash_0.x7.neg_mid VDPWR.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X78 flash_0.x4.VOUT flash_0.x4.VDPWR1 flash_0.x4.vintp flash_0.x7.VPRGPOS.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X79 flash_0.x3.stage2 flash_0.x3.stage1 flash_0.x3.stage1 flash_0.x3.stage1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X80 flash_0.x2.clkinb clk.t2 VAPWR.t1 VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X81 flash_0.x4.VOUT flash_0.x4.neg_mid_b.t14 flash_0.x4.dcgint.t4 flash_0.x4.dcgint.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X82 flash_0.x7.neg_mid_b.t6 flash_0.x7.neg_mid flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=1
X83 flash_0.x4.vintp flash_0.x4.pos_mid_b.t5 flash_0.x7.VPRGPOS.t20 flash_0.x7.VPRGPOS.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X84 VGND.t69 flash_0.x7.pos_en_b.t5 flash_0.x7.pos_mid VGND.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X85 flash_0.x7.dcgint.t7 flash_0.x7.neg_mid_b.t8 flash_0.x7.VOUT.t10 flash_0.x7.dcgint.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X86 flash_0.x3.clkb.t0 flash_0.x3.clkinb VAPWR.t12 VAPWR.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X87 flash_0.x7.vintp flash_0.x7.VDPWR1 flash_0.x7.VOUT.t5 flash_0.x7.VPRGPOS.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X88 flash_0.x7.VOUT.t8 VDPWR.t60 a_20416_28577# flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X89 flash_0.x4.vintp flash_0.x4.VDPWR1 flash_0.x4.VOUT flash_0.x7.VPRGPOS.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X90 flash_0.x7.VPRGPOS.t9 flash_0.x4.pos_mid_b.t6 flash_0.x4.vintp flash_0.x7.VPRGPOS.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X91 flash_0.x2.clkb flash_0.x2.stage2 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X92 flash_0.x2.stage1 flash_0.x2.stage1 VGND.t16 flash_0.x2.stage1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X93 flash_0.x7.VPRGPOS.t10 flash_0.x3.stage2 flash_0.x3.stage2 flash_0.x3.stage2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X94 VGND.t68 flash_0.x7.pos_en_b.t5 flash_0.x7.pos_mid VGND.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X95 flash_0.x4.pos_mid_b.t2 ui_in[0].t11 VGND.t61 VGND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X96 flash_0.x4.pos_mid flash_0.x4.pos_en_b.t5 VGND.t3 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X97 flash_0.x2.clkb.t1 flash_0.x2.clkinb VGND.t44 VGND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X98 flash_0.x3.clkina flash_0.x3.clkinb VAPWR.t10 VAPWR.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X99 flash_0.x7.vintp flash_0.x7.pos_mid_b.t8 flash_0.x7.VPRGPOS.t26 flash_0.x7.VPRGPOS.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X100 VDPWR.t46 flash_0.x4.neg_en_b.t8 flash_0.x4.neg_mid_b.t3 VDPWR.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X101 flash_0.x7.VOUT.t7 VDPWR.t61 a_20416_28577# flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X102 flash_0.x4.vintp flash_0.x4.pos_mid_b.t7 flash_0.x7.VPRGPOS.t7 flash_0.x7.VPRGPOS.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X103 flash_0.x7.dcgint.t11 flash_0.x7.pos_en_b.t6 VGND.t32 VGND.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X104 a_20416_28577# flash_0.x7.neg_mid_b.t9 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X105 flash_0.x2.clka.t0 flash_0.x2.clkina VAPWR.t13 VAPWR.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
X106 VGND.t34 ui_in[0].t12 flash_0.x7.neg_en_b.t1 VGND.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X107 flash_0.x7.neg_mid_b.t2 flash_0.x7.neg_en_b.t7 VDPWR.t14 VDPWR.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X108 flash_0.x4.pos_mid_b.t1 ui_in[0].t13 VGND.t35 VGND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X109 flash_0.x4.neg_mid ui_in[1].t12 VDPWR.t33 VDPWR.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X110 flash_0.x4.pos_mid flash_0.x4.pos_en_b.t5 VGND.t2 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X111 VDPWR.t31 ui_in[1].t13 flash_0.x4.neg_mid VDPWR.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X112 flash_0.x2.clka flash_0.x2.stage1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X113 flash_0.x7.VPRGPOS VGND.t37 sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X114 VDPWR.t45 flash_0.x4.neg_en_b.t9 flash_0.x4.neg_mid_b.t1 VDPWR.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X115 flash_0.x7.dcgint.t10 flash_0.x7.pos_en_b.t6 VGND.t30 VGND.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X116 a_20416_28577# flash_0.x7.neg_mid_b.t10 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X117 flash_0.x7.VOUT.t12 flash_0.x7.neg_mid_b.t11 flash_0.x7.dcgint.t5 flash_0.x7.dcgint.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X118 VDPWR.t1 ui_in[0].t14 flash_0.x7.neg_mid VDPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X119 flash_0.x7.neg_mid_b.t1 flash_0.x7.neg_en_b.t8 VDPWR.t16 VDPWR.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X120 flash_0.x4.neg_en_b.t2 ui_in[1].t14 VGND.t26 VGND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X121 flash_0.x4.pos_en_b.t2 ui_in[0].t15 VGND.t1 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X122 flash_0.x4.neg_mid ui_in[1].t15 VDPWR.t29 VDPWR.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X123 VDPWR.t54 ui_in[0].t16 flash_0.x7.neg_en_b.t3 VDPWR.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X124 flash_0.x7.dcgint.t4 flash_0.x7.neg_mid_b.t12 flash_0.x7.VOUT.t13 flash_0.x7.dcgint.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X125 flash_0.x2.clkinb clk.t3 VGND.t18 VGND.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X126 flash_0.x7.VOUT.t14 flash_0.x7.neg_mid_b.t13 flash_0.x7.dcgint.t3 flash_0.x7.dcgint.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X127 flash_0.x4.VOUT flash_0.x4.VDPWR1 flash_0.x4.vintp flash_0.x7.VPRGPOS.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X128 flash_0.x7.dcgint.t9 flash_0.x7.pos_en_b.t6 VGND.t28 VGND.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X129 flash_0.x3.clka.t1 flash_0.x3.clkina VGND.t65 VGND.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X130 flash_0.x5.A.t2 flash_0.x5.A.t0 a_9352_28387# flash_0.x5.A.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.5
X131 flash_0.x7.dcgint.t1 flash_0.x7.neg_mid_b.t14 flash_0.x7.VOUT.t9 flash_0.x7.dcgint.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X132 flash_0.x7.neg_mid_b.t0 flash_0.x7.neg_en_b.t9 VDPWR.t10 VDPWR.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X133 flash_0.x7.vintp flash_0.x7.VDPWR1 flash_0.x7.VOUT.t4 flash_0.x7.VPRGPOS.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X134 flash_0.x4.neg_en_b.t1 ui_in[1].t16 VDPWR.t27 VDPWR.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=3
X135 flash_0.x4.pos_en_b.t0 ui_in[0].t17 VDPWR.t23 VDPWR.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X136 VGND.t67 flash_0.x4.pos_en_b.t6 flash_0.x4.pos_mid VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X137 flash_0.x7.VPRGNEG flash_0.x7.neg_mid_b.t15 flash_0.x7.neg_mid flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.145 ps=1.58 w=0.5 l=1
X138 flash_0.x7.VOUT.t3 flash_0.x7.VDPWR1 flash_0.x7.vintp flash_0.x7.VPRGPOS.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X139 flash_0.x2.stage2 flash_0.x2.stage2 flash_0.x2.stage1 flash_0.x2.stage2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X140 flash_0.x7.VPRGPOS.t18 flash_0.x4.pos_mid_b.t8 flash_0.x4.vintp flash_0.x7.VPRGPOS.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X141 flash_0.x4.neg_mid ui_in[1].t17 VDPWR.t25 VDPWR.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X142 flash_0.x7.vintp flash_0.x7.pos_mid_b.t9 flash_0.x7.VPRGPOS.t25 flash_0.x7.VPRGPOS.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X143 flash_0.x7.VOUT.t2 flash_0.x7.VDPWR1 flash_0.x7.vintp flash_0.x7.VPRGPOS.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X144 flash_0.x7.VPRGPOS.t24 flash_0.x7.pos_mid_b flash_0.x7.pos_mid flash_0.x7.VPRGPOS.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X145 flash_0.x7.VPRGPOS.t31 flash_0.x4.pos_mid_b flash_0.x4.pos_mid flash_0.x7.VPRGPOS.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X146 VGND.t66 flash_0.x4.pos_en_b.t6 flash_0.x4.pos_mid VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X147 uo_out[0].t1 flash_0.x5.A.t5 VGND.t23 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X148 flash_0.x3.clkina flash_0.x3.clkinb VGND.t48 VGND.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X149 flash_0.x7.vintp flash_0.x7.VDPWR1 flash_0.x7.VOUT.t1 flash_0.x7.VPRGPOS.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X150 flash_0.x7.VPRGPOS.t22 flash_0.x7.pos_mid_b.t10 flash_0.x7.vintp flash_0.x7.VPRGPOS.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X151 flash_0.x6.Y.t0 ui_in[2].t2 VDPWR.t12 VDPWR.t11 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X152 flash_0.x7.VPRGNEG flash_0.x7.VPRGNEG flash_0.x2.stage2 flash_0.x7.VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
R0 VGND.t53 VGND.n121 1.77808e+07
R1 VGND.n205 VGND.n204 1.32662e+07
R2 VGND.n121 VGND.t27 9.06413e+06
R3 VGND.n205 VGND.n24 7.77048e+06
R4 VGND.n138 VGND.n129 136400
R5 VGND.n149 VGND.n118 77206.1
R6 VGND.n172 VGND.n63 55379.3
R7 VGND.n140 VGND.n139 41452.9
R8 VGND.n136 VGND.n135 28158.7
R9 VGND.n82 VGND.n67 26564
R10 VGND.n143 VGND.n129 26182
R11 VGND.n82 VGND.n81 19464
R12 VGND.n139 VGND.n138 18707.2
R13 VGND.n171 VGND.n170 17794
R14 VGND.n206 VGND.n22 17579
R15 VGND.n45 VGND.n41 17010.2
R16 VGND.n52 VGND.n41 17010.2
R17 VGND.n183 VGND.n56 17010.2
R18 VGND.n174 VGND.n56 17010.2
R19 VGND.n145 VGND.n129 16052.9
R20 VGND.n136 VGND.n22 15944.1
R21 VGND.n170 VGND.n82 15655.2
R22 VGND.n152 VGND.n118 15267.5
R23 VGND.n172 VGND.n171 13983.9
R24 VGND.n171 VGND.n64 12678.4
R25 VGND.n138 VGND.n137 11203.8
R26 VGND.n207 VGND.n206 8682.25
R27 VGND.n152 VGND.n151 8288.46
R28 VGND.n71 VGND.n22 7672.91
R29 VGND.n128 VGND.t57 6465.71
R30 VGND.n137 VGND.n118 5878.85
R31 VGND.n205 VGND.n23 5801.34
R32 VGND.n58 VGND.n55 5607.68
R33 VGND.n43 VGND.n40 5607.68
R34 VGND.n40 VGND.n23 5607.68
R35 VGND.n62 VGND.n55 5607.68
R36 VGND.n120 VGND.n119 5067.26
R37 VGND.n141 VGND.n140 4557.14
R38 VGND.t33 VGND.t6 4288.33
R39 VGND.t6 VGND.t14 4288.33
R40 VGND.t4 VGND.t0 4288.33
R41 VGND.t0 VGND.t9 4288.33
R42 VGND.n168 VGND.n83 3957.38
R43 VGND.n168 VGND.n84 3957.38
R44 VGND.n133 VGND.n84 3957.38
R45 VGND.n133 VGND.n83 3957.38
R46 VGND.n72 VGND.n68 3957.38
R47 VGND.n72 VGND.n69 3957.38
R48 VGND.n80 VGND.n69 3957.38
R49 VGND.n80 VGND.n68 3957.38
R50 VGND.n203 VGND.n25 3790.36
R51 VGND.n60 VGND.n25 3790.36
R52 VGND.n189 VGND.n188 3790.36
R53 VGND.n188 VGND.n38 3790.36
R54 VGND.n148 VGND.t12 3495.43
R55 VGND.n142 VGND.t25 3495.43
R56 VGND.n81 VGND.t62 3200.66
R57 VGND.n71 VGND.t62 3200.66
R58 VGND.n149 VGND.n148 2827
R59 VGND.n143 VGND.n142 2827
R60 VGND.n43 VGND.n39 2736.73
R61 VGND.n147 VGND.n145 2648.22
R62 VGND.n139 VGND.n135 2546
R63 VGND.t14 VGND.n147 2345.18
R64 VGND.t9 VGND.n141 2345.18
R65 VGND.n172 VGND.n62 2341.85
R66 VGND.n151 VGND.t12 2331.85
R67 VGND.n63 VGND.n58 2309.11
R68 VGND.n54 VGND.n53 2233.78
R69 VGND.n137 VGND.n136 2176.84
R70 VGND.n206 VGND.n205 1977.24
R71 VGND.n208 VGND.n20 1900.12
R72 VGND.n208 VGND.n21 1900.12
R73 VGND.n66 VGND.n21 1900.12
R74 VGND.n66 VGND.n20 1900.12
R75 VGND.n185 VGND.n184 1830.35
R76 VGND.t25 VGND.n128 1820.3
R77 VGND.n140 VGND.n64 1788.04
R78 VGND.n135 VGND.n134 1768.36
R79 VGND.n44 VGND.n23 1501.04
R80 VGND.n54 VGND.n39 1195.35
R81 VGND.n170 VGND.n169 1151.51
R82 VGND.n51 VGND.n42 1139.95
R83 VGND.n46 VGND.n42 1139.95
R84 VGND.n182 VGND.n57 1139.95
R85 VGND.n175 VGND.n57 1139.95
R86 VGND.t31 VGND.n152 1094.37
R87 VGND.n134 VGND.t22 1089.55
R88 VGND.n169 VGND.t22 1089.55
R89 VGND.n120 VGND.n54 931.699
R90 VGND.n62 VGND.n61 883.615
R91 VGND.n148 VGND.t33 792.894
R92 VGND.n142 VGND.t4 792.894
R93 VGND.t43 VGND.t51 757.616
R94 VGND.n67 VGND.t59 660
R95 VGND.n207 VGND.t59 660
R96 VGND.n173 VGND.n58 657.409
R97 VGND.n15 VGND.t41 650.87
R98 VGND.t45 VGND.t17 597.753
R99 VGND.n121 VGND.n120 522.082
R100 VGND.t57 VGND.t55 487.856
R101 VGND.n61 VGND.t43 478.974
R102 VGND.t64 VGND.t49 470.42
R103 VGND.n202 VGND.n201 437.836
R104 VGND.n201 VGND.n27 437.836
R105 VGND.n191 VGND.n37 437.836
R106 VGND.n191 VGND.n190 437.836
R107 VGND.n204 VGND.t17 424.973
R108 VGND.n44 VGND.n43 417.728
R109 VGND.n185 VGND.n54 402.44
R110 VGND.t51 VGND.n59 378.808
R111 VGND.n59 VGND.t45 378.808
R112 VGND.t47 VGND.t20 350.719
R113 VGND.n127 VGND.t53 304.329
R114 VGND.t49 VGND.n186 297.404
R115 VGND.n132 VGND.n131 257.13
R116 VGND.n132 VGND.n86 257.13
R117 VGND.n79 VGND.n70 257.13
R118 VGND.n79 VGND.n78 257.13
R119 VGND.n187 VGND.t64 235.209
R120 VGND.n157 VGND.t28 230.898
R121 VGND.n155 VGND.t30 230.898
R122 VGND.n156 VGND.t32 230.898
R123 VGND.n125 VGND.t54 230.898
R124 VGND.n122 VGND.t56 230.898
R125 VGND.n123 VGND.t58 230.898
R126 VGND.n131 VGND.n85 229.272
R127 VGND.n166 VGND.n86 229.272
R128 VGND.n74 VGND.n70 229.272
R129 VGND.n78 VGND.n77 229.272
R130 VGND.n193 VGND.t48 227.643
R131 VGND.n199 VGND.t46 227.643
R132 VGND.n26 VGND.t18 227.398
R133 VGND.n34 VGND.t21 227.398
R134 VGND.n187 VGND.t47 222.901
R135 VGND.n209 VGND.n19 221.742
R136 VGND.n65 VGND.n19 221.742
R137 VGND.n65 VGND.n18 221.742
R138 VGND.t20 VGND.n24 221.728
R139 VGND.n144 VGND.n143 193.178
R140 VGND.n150 VGND.n149 193.178
R141 VGND.t55 VGND.n127 183.528
R142 VGND.n145 VGND.n144 182.445
R143 VGND.n151 VGND.n150 182.445
R144 VGND.t29 VGND.t31 157.787
R145 VGND.n210 VGND.n18 152.194
R146 VGND.n147 VGND.n146 152.111
R147 VGND.n141 VGND.n130 152.111
R148 VGND.n135 VGND.n64 147.569
R149 VGND.n20 VGND.n18 146.25
R150 VGND.t59 VGND.n20 146.25
R151 VGND.n21 VGND.n19 146.25
R152 VGND.t59 VGND.n21 146.25
R153 VGND.n133 VGND.n132 117.001
R154 VGND.n134 VGND.n133 117.001
R155 VGND.n168 VGND.n167 117.001
R156 VGND.n169 VGND.n168 117.001
R157 VGND.n80 VGND.n79 117.001
R158 VGND.n81 VGND.n80 117.001
R159 VGND.n73 VGND.n72 117.001
R160 VGND.n72 VGND.n71 117.001
R161 VGND.n186 VGND.n185 107.427
R162 VGND.n53 VGND.n40 102.35
R163 VGND.n184 VGND.n55 102.35
R164 VGND.n153 VGND.t27 98.4295
R165 VGND.n60 VGND.n27 97.5005
R166 VGND.n61 VGND.n60 97.5005
R167 VGND.n203 VGND.n202 97.5005
R168 VGND.n204 VGND.n203 97.5005
R169 VGND.n38 VGND.n37 97.5005
R170 VGND.n186 VGND.n38 97.5005
R171 VGND.n190 VGND.n189 97.5005
R172 VGND.n189 VGND.n24 97.5005
R173 VGND.n115 VGND.n114 97.1505
R174 VGND.n108 VGND.n107 97.1505
R175 VGND.n111 VGND.n110 97.1505
R176 VGND.n104 VGND.n103 97.1505
R177 VGND.n113 VGND.n112 97.1505
R178 VGND.n106 VGND.n105 97.1505
R179 VGND.n99 VGND.n98 97.1505
R180 VGND.n92 VGND.n91 97.1505
R181 VGND.n95 VGND.n94 97.1505
R182 VGND.n88 VGND.n87 97.1505
R183 VGND.n97 VGND.n96 97.1505
R184 VGND.n90 VGND.n89 97.1505
R185 VGND.n119 VGND.n63 95.855
R186 VGND.n114 VGND.t19 95.7605
R187 VGND.n114 VGND.t24 95.7605
R188 VGND.n107 VGND.t39 95.7605
R189 VGND.n107 VGND.t34 95.7605
R190 VGND.n110 VGND.t7 95.7605
R191 VGND.n110 VGND.t70 95.7605
R192 VGND.n103 VGND.t36 95.7605
R193 VGND.n103 VGND.t68 95.7605
R194 VGND.n112 VGND.t8 95.7605
R195 VGND.n112 VGND.t15 95.7605
R196 VGND.n105 VGND.t13 95.7605
R197 VGND.n105 VGND.t69 95.7605
R198 VGND.n98 VGND.t1 95.7605
R199 VGND.n98 VGND.t38 95.7605
R200 VGND.n91 VGND.t26 95.7605
R201 VGND.n91 VGND.t5 95.7605
R202 VGND.n94 VGND.t2 95.7605
R203 VGND.n94 VGND.t10 95.7605
R204 VGND.n87 VGND.t35 95.7605
R205 VGND.n87 VGND.t66 95.7605
R206 VGND.n96 VGND.t3 95.7605
R207 VGND.n96 VGND.t11 95.7605
R208 VGND.n89 VGND.t61 95.7605
R209 VGND.n89 VGND.t67 95.7605
R210 VGND.n164 VGND.t23 83.754
R211 VGND.n76 VGND.t63 83.7172
R212 VGND.n36 VGND.t50 83.1807
R213 VGND.n28 VGND.t44 83.1807
R214 VGND.n35 VGND.t65 82.9558
R215 VGND.n29 VGND.t52 82.9558
R216 VGND.n30 VGND.t16 82.8472
R217 VGND.n154 VGND.n153 73.7068
R218 VGND.n127 VGND.n126 73.7068
R219 VGND.n66 VGND.n65 65.0005
R220 VGND.n67 VGND.n66 65.0005
R221 VGND.n209 VGND.n208 65.0005
R222 VGND.n208 VGND.n207 65.0005
R223 VGND.n153 VGND.t29 59.3584
R224 VGND.n210 VGND.n209 56.9466
R225 VGND.n131 VGND.n83 53.1823
R226 VGND.n83 VGND.t22 53.1823
R227 VGND.n86 VGND.n84 53.1823
R228 VGND.n84 VGND.t22 53.1823
R229 VGND.n70 VGND.n68 53.1823
R230 VGND.n68 VGND.t62 53.1823
R231 VGND.n78 VGND.n69 53.1823
R232 VGND.n69 VGND.t62 53.1823
R233 VGND.n211 VGND.t60 41.2645
R234 VGND.n167 VGND.n85 27.8593
R235 VGND.n167 VGND.n166 27.8593
R236 VGND.n74 VGND.n73 27.8593
R237 VGND.n77 VGND.n73 27.8593
R238 VGND.n57 VGND.n56 26.5914
R239 VGND.n119 VGND.n56 26.5914
R240 VGND.n42 VGND.n41 26.5914
R241 VGND.n41 VGND.n39 26.5914
R242 VGND.n201 VGND.n25 24.3755
R243 VGND.n59 VGND.n25 24.3755
R244 VGND.n191 VGND.n188 24.3755
R245 VGND.n188 VGND.n187 24.3755
R246 VGND.n173 VGND.n172 20.4593
R247 VGND.n75 VGND.n74 9.35514
R248 VGND.n77 VGND 9.33194
R249 VGND.n166 VGND.n165 9.3005
R250 VGND.n165 VGND.n85 9.3005
R251 VGND.n46 VGND.n45 9.28621
R252 VGND.n45 VGND.n44 9.28621
R253 VGND.n183 VGND.n182 9.28621
R254 VGND.n184 VGND.n183 9.28621
R255 VGND.n52 VGND.n51 9.28621
R256 VGND.n53 VGND.n52 9.28621
R257 VGND.n175 VGND.n174 9.28621
R258 VGND.n174 VGND.n173 9.28621
R259 VGND.n213 VGND.n16 8.39735
R260 VGND.n48 VGND.n47 8.21246
R261 VGND.n181 VGND.n180 8.21246
R262 VGND.n49 VGND.n48 7.33652
R263 VGND.n180 VGND.n179 7.33652
R264 VGND.n146 VGND.n117 6.24424
R265 VGND.n130 VGND.n101 6.24424
R266 VGND.n47 VGND 5.82387
R267 VGND.n181 VGND 5.82387
R268 VGND.n212 VGND.n211 5.18907
R269 VGND.n50 VGND 5.15194
R270 VGND.n176 VGND 5.15194
R271 VGND.n164 VGND.n163 5.15155
R272 VGND.n15 VGND.t40 4.756
R273 VGND.n124 VGND.n123 4.5005
R274 VGND.n124 VGND.n122 4.5005
R275 VGND.n125 VGND.n124 4.5005
R276 VGND.n158 VGND.n156 4.5005
R277 VGND.n158 VGND.n155 4.5005
R278 VGND.n158 VGND.n157 4.5005
R279 VGND.n33 VGND.n32 4.12801
R280 VGND.n178 VGND.n177 4.12801
R281 VGND.n147 VGND.n128 4.11265
R282 VGND.n196 VGND 3.81988
R283 VGND.n215 VGND 3.32011
R284 VGND.n37 VGND.n36 3.31952
R285 VGND.n28 VGND.n27 3.31952
R286 VGND.n195 VGND.n33 3.218
R287 VGND.n16 VGND.n15 3.20171
R288 VGND.n160 VGND.n159 3.12737
R289 VGND.n162 VGND.n161 3.00925
R290 uio_oe[7] VGND.n215 2.60868
R291 VGND.n211 VGND.n210 2.3255
R292 VGND.n109 VGND.n106 2.2505
R293 VGND.n116 VGND.n113 2.2505
R294 VGND.n109 VGND.n104 2.2505
R295 VGND.n116 VGND.n111 2.2505
R296 VGND.n109 VGND.n108 2.2505
R297 VGND.n116 VGND.n115 2.2505
R298 VGND.n93 VGND.n90 2.2505
R299 VGND.n100 VGND.n97 2.2505
R300 VGND.n93 VGND.n88 2.2505
R301 VGND.n100 VGND.n95 2.2505
R302 VGND.n93 VGND.n92 2.2505
R303 VGND.n100 VGND.n99 2.2505
R304 VGND.n126 VGND.n125 2.04916
R305 VGND.n157 VGND.n154 2.04916
R306 VGND.n163 VGND.n162 2.00487
R307 VGND.n178 VGND.n31 1.913
R308 VGND.n163 VGND.n17 1.74613
R309 VGND.n31 VGND.n30 1.5555
R310 VGND.n202 VGND.n26 1.5505
R311 VGND.n190 VGND.n34 1.5505
R312 VGND.n160 VGND.n117 1.31425
R313 VGND.n197 VGND.n31 1.3055
R314 VGND.n162 VGND.n101 1.248
R315 VGND.n212 VGND.n17 1.188
R316 VGND.n196 VGND.n17 1.1555
R317 VGND.n36 VGND.n35 0.879043
R318 VGND.n29 VGND.n28 0.879043
R319 VGND.n215 VGND.n214 0.751794
R320 VGND.n213 VGND.n212 0.525188
R321 VGND.n198 VGND.n197 0.501003
R322 VGND.n195 VGND.n194 0.501003
R323 VGND.n48 VGND.n42 0.443357
R324 VGND.n180 VGND.n57 0.443357
R325 VGND.n201 VGND.n200 0.404848
R326 VGND.n192 VGND.n191 0.404848
R327 VGND.n116 VGND.n109 0.378453
R328 VGND.n100 VGND.n93 0.378453
R329 VGND.n159 VGND.n154 0.285933
R330 VGND.n126 VGND.n102 0.28175
R331 VGND.n161 VGND.n160 0.27425
R332 VGND.n161 VGND.n102 0.236484
R333 VGND.n200 VGND.n199 0.221088
R334 VGND.n193 VGND.n192 0.221088
R335 VGND.n199 VGND 0.214961
R336 VGND VGND.n193 0.214961
R337 VGND.n124 VGND 0.204732
R338 VGND VGND.n158 0.204732
R339 VGND VGND.n196 0.177375
R340 VGND.n75 VGND.n16 0.168469
R341 VGND.n214 VGND.n213 0.166437
R342 VGND.n0 uo_out[1] 0.16627
R343 VGND.n1 uo_out[2] 0.16627
R344 VGND.n2 uo_out[3] 0.16627
R345 VGND.n3 uo_out[4] 0.16627
R346 VGND.n4 uo_out[5] 0.16627
R347 VGND.n5 uo_out[6] 0.16627
R348 VGND.n6 uo_out[7] 0.16627
R349 VGND.n7 uio_out[0] 0.16627
R350 VGND.n8 uio_out[1] 0.16627
R351 VGND.n9 uio_out[2] 0.16627
R352 VGND.n10 uio_out[3] 0.16627
R353 VGND.n11 uio_out[4] 0.16627
R354 VGND.n12 uio_out[5] 0.16627
R355 VGND.n13 uio_out[6] 0.16627
R356 VGND.n14 uio_out[7] 0.16627
R357 uio_oe[0] VGND.n222 0.16627
R358 uio_oe[1] VGND.n221 0.16627
R359 uio_oe[2] VGND.n220 0.16627
R360 uio_oe[3] VGND.n219 0.16627
R361 uio_oe[4] VGND.n218 0.16627
R362 uio_oe[5] VGND.n217 0.16627
R363 uio_oe[6] VGND.n216 0.16627
R364 VGND.n146 VGND 0.157483
R365 VGND.n130 VGND 0.157483
R366 VGND.n50 VGND.n49 0.15675
R367 VGND.n179 VGND.n176 0.15675
R368 VGND.n47 VGND.n46 0.1555
R369 VGND.n51 VGND.n50 0.1555
R370 VGND.n182 VGND.n181 0.1555
R371 VGND.n176 VGND.n175 0.1555
R372 VGND.n115 VGND 0.102773
R373 VGND.n108 VGND 0.102773
R374 VGND.n111 VGND 0.102773
R375 VGND.n104 VGND 0.102773
R376 VGND.n113 VGND 0.102773
R377 VGND.n106 VGND 0.102773
R378 VGND.n99 VGND 0.102773
R379 VGND.n92 VGND 0.102773
R380 VGND.n95 VGND 0.102773
R381 VGND.n88 VGND 0.102773
R382 VGND.n97 VGND 0.102773
R383 VGND.n90 VGND 0.102773
R384 VGND.n198 VGND.n26 0.0904491
R385 VGND.n194 VGND.n34 0.0904491
R386 VGND VGND.n198 0.0659475
R387 VGND.n194 VGND 0.0659475
R388 VGND.n49 VGND.n33 0.0657174
R389 VGND.n179 VGND.n178 0.0657174
R390 VGND.n214 VGND 0.062375
R391 VGND.n30 VGND 0.0609396
R392 VGND VGND.n195 0.05925
R393 VGND.n197 VGND 0.05925
R394 VGND.n155 VGND 0.0544773
R395 VGND.n156 VGND 0.0544773
R396 VGND.n122 VGND 0.0544773
R397 VGND.n123 VGND 0.0544773
R398 VGND.n125 VGND 0.048
R399 VGND.n157 VGND 0.048
R400 VGND.n165 VGND.n164 0.034875
R401 VGND.n177 VGND.t42 0.0314016
R402 VGND.n32 VGND.t37 0.0314016
R403 VGND VGND.n102 0.0312579
R404 VGND.n0 uo_out[2] 0.0302667
R405 VGND.n1 uo_out[3] 0.0302667
R406 VGND.n2 uo_out[4] 0.0302667
R407 VGND.n3 uo_out[5] 0.0302667
R408 VGND.n4 uo_out[6] 0.0302667
R409 VGND.n5 uo_out[7] 0.0302667
R410 VGND.n6 uio_out[0] 0.0302667
R411 VGND.n7 uio_out[1] 0.0302667
R412 VGND.n8 uio_out[2] 0.0302667
R413 VGND.n9 uio_out[3] 0.0302667
R414 VGND.n10 uio_out[4] 0.0302667
R415 VGND.n11 uio_out[5] 0.0302667
R416 VGND.n12 uio_out[6] 0.0302667
R417 VGND.n13 uio_out[7] 0.0302667
R418 VGND.n14 uio_oe[0] 0.0302667
R419 VGND.n222 uio_oe[1] 0.0302667
R420 VGND.n221 uio_oe[2] 0.0302667
R421 VGND.n220 uio_oe[3] 0.0302667
R422 VGND.n219 uio_oe[4] 0.0302667
R423 VGND.n218 uio_oe[5] 0.0302667
R424 VGND.n217 uio_oe[6] 0.0302667
R425 VGND.n216 uio_oe[7] 0.0302667
R426 VGND.n159 VGND 0.0270748
R427 VGND VGND.n76 0.0244521
R428 VGND.n150 VGND 0.0234785
R429 VGND.n144 VGND 0.0234785
R430 VGND.n200 VGND.n29 0.0194951
R431 VGND.n192 VGND.n35 0.0194951
R432 VGND.n117 VGND.n116 0.0182165
R433 VGND.n101 VGND.n100 0.0182165
R434 uo_out[2] VGND.n0 0.010027
R435 uo_out[3] VGND.n1 0.010027
R436 uo_out[4] VGND.n2 0.010027
R437 uo_out[5] VGND.n3 0.010027
R438 uo_out[6] VGND.n4 0.010027
R439 uo_out[7] VGND.n5 0.010027
R440 uio_out[0] VGND.n6 0.010027
R441 uio_out[1] VGND.n7 0.010027
R442 uio_out[2] VGND.n8 0.010027
R443 uio_out[3] VGND.n9 0.010027
R444 uio_out[4] VGND.n10 0.010027
R445 uio_out[5] VGND.n11 0.010027
R446 uio_out[6] VGND.n12 0.010027
R447 uio_out[7] VGND.n13 0.010027
R448 uio_oe[0] VGND.n14 0.010027
R449 VGND.n222 uio_oe[1] 0.010027
R450 VGND.n221 uio_oe[2] 0.010027
R451 VGND.n220 uio_oe[3] 0.010027
R452 VGND.n219 uio_oe[4] 0.010027
R453 VGND.n218 uio_oe[5] 0.010027
R454 VGND.n217 uio_oe[6] 0.010027
R455 VGND.n216 uio_oe[7] 0.010027
R456 VGND.n165 VGND 0.008625
R457 VGND.n76 VGND.n75 0.0012485
R458 VGND.n177 VGND 0.000981102
R459 VGND.n32 VGND 0.000981102
R460 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t3 649.691
R461 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t2 227.442
R462 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t4 227.442
R463 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t1 227.361
R464 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t0 227.361
R465 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t9 216.731
R466 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t10 216.731
R467 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t8 216.731
R468 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t5 216.731
R469 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t6 216.731
R470 flash_0.x7.pos_mid_b flash_0.x7.pos_mid_b.t7 216.731
R471 flash_0.x7.VPRGPOS.n6 flash_0.x7.VPRGPOS.n4 4689.72
R472 flash_0.x7.VPRGPOS.n9 flash_0.x7.VPRGPOS.n8 4689.72
R473 flash_0.x7.VPRGPOS.n7 flash_0.x7.VPRGPOS.n6 1828.1
R474 flash_0.x7.VPRGPOS.n9 flash_0.x7.VPRGPOS.n3 1828.1
R475 flash_0.x7.VPRGPOS.n5 flash_0.x7.VPRGPOS.n1 902.777
R476 flash_0.x7.VPRGPOS.n5 flash_0.x7.VPRGPOS.n2 902.777
R477 flash_0.x7.VPRGPOS.n10 flash_0.x7.VPRGPOS.n2 880.232
R478 flash_0.x7.VPRGPOS.n11 flash_0.x7.VPRGPOS.n1 874.658
R479 flash_0.x7.VPRGPOS.t14 flash_0.x7.VPRGPOS.t23 809.375
R480 flash_0.x7.VPRGPOS.t19 flash_0.x7.VPRGPOS.t2 809.375
R481 flash_0.x7.VPRGPOS.n12 flash_0.x7.VPRGPOS.t1 649.856
R482 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t18 649.715
R483 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t27 649.715
R484 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t30 649.691
R485 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t24 649.691
R486 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t3 649.691
R487 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t31 649.691
R488 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t20 649.691
R489 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t25 649.691
R490 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n14 594.301
R491 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n13 594.301
R492 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n18 594.301
R493 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n19 594.301
R494 flash_0.x7.VPRGPOS.t11 flash_0.x7.VPRGPOS.t16 246.875
R495 flash_0.x7.VPRGPOS.t12 flash_0.x7.VPRGPOS.t11 246.875
R496 flash_0.x7.VPRGPOS.t15 flash_0.x7.VPRGPOS.t12 246.875
R497 flash_0.x7.VPRGPOS.t13 flash_0.x7.VPRGPOS.t15 246.875
R498 flash_0.x7.VPRGPOS.t6 flash_0.x7.VPRGPOS.t17 246.875
R499 flash_0.x7.VPRGPOS.t4 flash_0.x7.VPRGPOS.t6 246.875
R500 flash_0.x7.VPRGPOS.t21 flash_0.x7.VPRGPOS.t4 246.875
R501 flash_0.x7.VPRGPOS.t8 flash_0.x7.VPRGPOS.t21 246.875
R502 flash_0.x7.VPRGPOS.n0 flash_0.x7.VPRGPOS.t13 237.5
R503 flash_0.x7.VPRGPOS.n15 flash_0.x7.VPRGPOS.t8 237.5
R504 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.t10 82.8472
R505 flash_0.x7.VPRGPOS.n14 flash_0.x7.VPRGPOS.t32 55.3905
R506 flash_0.x7.VPRGPOS.n14 flash_0.x7.VPRGPOS.t9 55.3905
R507 flash_0.x7.VPRGPOS.n13 flash_0.x7.VPRGPOS.t7 55.3905
R508 flash_0.x7.VPRGPOS.n13 flash_0.x7.VPRGPOS.t5 55.3905
R509 flash_0.x7.VPRGPOS.n18 flash_0.x7.VPRGPOS.t26 55.3905
R510 flash_0.x7.VPRGPOS.n18 flash_0.x7.VPRGPOS.t22 55.3905
R511 flash_0.x7.VPRGPOS.n19 flash_0.x7.VPRGPOS.t28 55.3905
R512 flash_0.x7.VPRGPOS.n19 flash_0.x7.VPRGPOS.t29 55.3905
R513 flash_0.x7.VPRGPOS.n6 flash_0.x7.VPRGPOS.n5 37.0005
R514 flash_0.x7.VPRGPOS.n10 flash_0.x7.VPRGPOS.n9 37.0005
R515 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n0 16.1367
R516 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n15 16.1367
R517 flash_0.x7.VPRGPOS.n17 flash_0.x7.VPRGPOS 13.9898
R518 flash_0.x7.VPRGPOS.n0 flash_0.x7.VPRGPOS.t14 9.3755
R519 flash_0.x7.VPRGPOS.n15 flash_0.x7.VPRGPOS.t19 9.3755
R520 flash_0.x7.VPRGPOS.n4 flash_0.x7.VPRGPOS.n1 3.03329
R521 flash_0.x7.VPRGPOS.n8 flash_0.x7.VPRGPOS.n2 3.03329
R522 flash_0.x7.VPRGPOS.n16 flash_0.x7.VPRGPOS 2.77904
R523 flash_0.x7.VPRGPOS.n11 flash_0.x7.VPRGPOS.n10 2.70819
R524 flash_0.x7.VPRGPOS flash_0.x7.VPRGPOS.n17 2.54902
R525 flash_0.x7.VPRGPOS.n12 flash_0.x7.VPRGPOS.n11 1.8605
R526 flash_0.x7.VPRGPOS.n4 flash_0.x7.VPRGPOS.n3 1.85038
R527 flash_0.x7.VPRGPOS.n8 flash_0.x7.VPRGPOS.n7 1.85038
R528 flash_0.x7.VPRGPOS.n16 flash_0.x7.VPRGPOS.n12 1.79707
R529 flash_0.x7.VPRGPOS.n17 flash_0.x7.VPRGPOS.n16 1.40849
R530 flash_0.x7.VPRGPOS.t0 flash_0.x7.VPRGPOS.n3 1.18321
R531 flash_0.x7.VPRGPOS.n7 flash_0.x7.VPRGPOS.t0 1.18321
R532 VAPWR.n62 VAPWR.n4 2380.24
R533 VAPWR.n114 VAPWR.n73 2380.24
R534 VAPWR.n64 VAPWR.n4 2376.31
R535 VAPWR.n116 VAPWR.n73 2376.31
R536 VAPWR.n44 VAPWR.n42 2332.91
R537 VAPWR.n45 VAPWR.n44 2332.91
R538 VAPWR.n46 VAPWR.n45 2332.91
R539 VAPWR.n46 VAPWR.n42 2332.91
R540 VAPWR.n27 VAPWR.n25 2332.91
R541 VAPWR.n28 VAPWR.n27 2332.91
R542 VAPWR.n29 VAPWR.n28 2332.91
R543 VAPWR.n29 VAPWR.n25 2332.91
R544 VAPWR.n13 VAPWR.n12 2332.91
R545 VAPWR.n13 VAPWR.n11 2332.91
R546 VAPWR.n93 VAPWR.n92 2332.91
R547 VAPWR.n93 VAPWR.n91 2332.91
R548 VAPWR.n87 VAPWR.n83 1577.4
R549 VAPWR.n84 VAPWR.n81 1577.4
R550 VAPWR.n47 VAPWR.n38 1551.32
R551 VAPWR.n43 VAPWR.n38 1551.32
R552 VAPWR.n26 VAPWR.n24 1551.32
R553 VAPWR.n26 VAPWR.n21 1551.32
R554 VAPWR.n30 VAPWR.n21 1551.32
R555 VAPWR.n30 VAPWR.n24 1551.32
R556 VAPWR.n47 VAPWR.n41 1538.26
R557 VAPWR.n43 VAPWR.n41 1538.26
R558 VAPWR.n58 VAPWR.n7 1516.38
R559 VAPWR.n58 VAPWR.n6 1516.38
R560 VAPWR.n110 VAPWR.n76 1516.38
R561 VAPWR.n110 VAPWR.n75 1516.38
R562 VAPWR.n14 VAPWR.n7 1514.88
R563 VAPWR.n14 VAPWR.n6 1514.88
R564 VAPWR.n94 VAPWR.n76 1514.88
R565 VAPWR.n94 VAPWR.n75 1514.88
R566 VAPWR.n12 VAPWR.n5 1046.2
R567 VAPWR.n11 VAPWR.n5 1046.2
R568 VAPWR.n92 VAPWR.n74 1046.2
R569 VAPWR.n91 VAPWR.n74 1046.2
R570 VAPWR.n85 VAPWR.n84 722.497
R571 VAPWR.n87 VAPWR.n86 722.497
R572 VAPWR.n0 VAPWR.t6 649.99
R573 VAPWR.n121 VAPWR.t10 649.99
R574 VAPWR.n1 VAPWR.t1 649.765
R575 VAPWR.n71 VAPWR.t16 649.765
R576 VAPWR.t0 VAPWR.t5 487.901
R577 VAPWR.t15 VAPWR.t9 487.901
R578 VAPWR.n66 VAPWR.n3 460.425
R579 VAPWR.n118 VAPWR.n72 460.425
R580 VAPWR.n66 VAPWR.n65 459.671
R581 VAPWR.n118 VAPWR.n117 459.671
R582 VAPWR.n40 VAPWR.n37 386.635
R583 VAPWR.n48 VAPWR.n40 386.635
R584 VAPWR.n49 VAPWR.n37 386.635
R585 VAPWR.n23 VAPWR.n20 386.635
R586 VAPWR.n31 VAPWR.n23 386.635
R587 VAPWR.n32 VAPWR.n20 386.635
R588 VAPWR.n15 VAPWR.n8 386.635
R589 VAPWR.n15 VAPWR.n9 386.635
R590 VAPWR.n57 VAPWR.n8 386.635
R591 VAPWR.n57 VAPWR.n9 386.635
R592 VAPWR.n95 VAPWR.n77 386.635
R593 VAPWR.n95 VAPWR.n78 386.635
R594 VAPWR.n109 VAPWR.n78 386.635
R595 VAPWR.n109 VAPWR.n77 386.635
R596 VAPWR.n64 VAPWR.t0 331.582
R597 VAPWR.n116 VAPWR.t15 331.582
R598 VAPWR.n61 VAPWR.n60 251.28
R599 VAPWR.n113 VAPWR.n112 251.28
R600 VAPWR.t2 VAPWR 236.188
R601 VAPWR.n97 VAPWR.t2 236.011
R602 VAPWR.n49 VAPWR 195.012
R603 VAPWR.n32 VAPWR 195.012
R604 VAPWR VAPWR.n48 191.625
R605 VAPWR VAPWR.n31 191.625
R606 VAPWR.n106 VAPWR.n82 184.847
R607 VAPWR.n107 VAPWR.n106 184.847
R608 VAPWR.n107 VAPWR.n80 184.847
R609 VAPWR.n82 VAPWR.n80 184.847
R610 VAPWR.n59 VAPWR.n5 172.655
R611 VAPWR.n111 VAPWR.n74 172.655
R612 VAPWR.n55 VAPWR.t8 167.41
R613 VAPWR.n79 VAPWR.t12 167.41
R614 VAPWR.n120 VAPWR.t14 167.251
R615 VAPWR.n68 VAPWR.t13 167.141
R616 VAPWR.n60 VAPWR.n59 160.495
R617 VAPWR.n112 VAPWR.n111 160.495
R618 VAPWR.n107 VAPWR.n81 146.25
R619 VAPWR.n83 VAPWR.n82 146.25
R620 VAPWR.n106 VAPWR.n87 97.5005
R621 VAPWR.n84 VAPWR.n80 97.5005
R622 VAPWR.n105 VAPWR.t4 82.8472
R623 VAPWR.t5 VAPWR.t7 81.0585
R624 VAPWR.t9 VAPWR.t11 81.0585
R625 VAPWR.n85 VAPWR.n83 72.5386
R626 VAPWR.n86 VAPWR.n81 72.5386
R627 VAPWR.n86 VAPWR.t3 66.988
R628 VAPWR.t3 VAPWR.n85 66.988
R629 VAPWR.n63 VAPWR.n61 34.0449
R630 VAPWR.n115 VAPWR.n113 34.0449
R631 VAPWR.n62 VAPWR.n3 23.1255
R632 VAPWR.n63 VAPWR.n62 23.1255
R633 VAPWR.n65 VAPWR.n64 23.1255
R634 VAPWR.n114 VAPWR.n72 23.1255
R635 VAPWR.n115 VAPWR.n114 23.1255
R636 VAPWR.n117 VAPWR.n116 23.1255
R637 VAPWR.t5 VAPWR.n61 21.1116
R638 VAPWR.t9 VAPWR.n113 21.1116
R639 VAPWR.n43 VAPWR.n37 14.2313
R640 VAPWR.n44 VAPWR.n43 14.2313
R641 VAPWR.n48 VAPWR.n47 14.2313
R642 VAPWR.n47 VAPWR.n46 14.2313
R643 VAPWR.n26 VAPWR.n20 14.2313
R644 VAPWR.n27 VAPWR.n26 14.2313
R645 VAPWR.n31 VAPWR.n30 14.2313
R646 VAPWR.n30 VAPWR.n29 14.2313
R647 VAPWR.n15 VAPWR.n14 14.2313
R648 VAPWR.n14 VAPWR.n13 14.2313
R649 VAPWR.n58 VAPWR.n57 14.2313
R650 VAPWR.n59 VAPWR.n58 14.2313
R651 VAPWR.n95 VAPWR.n94 14.2313
R652 VAPWR.n94 VAPWR.n93 14.2313
R653 VAPWR.n110 VAPWR.n109 14.2313
R654 VAPWR.n111 VAPWR.n110 14.2313
R655 VAPWR.n41 VAPWR.n40 12.3338
R656 VAPWR.n42 VAPWR.n41 12.3338
R657 VAPWR.n49 VAPWR.n38 12.3338
R658 VAPWR.n45 VAPWR.n38 12.3338
R659 VAPWR.n24 VAPWR.n23 12.3338
R660 VAPWR.n25 VAPWR.n24 12.3338
R661 VAPWR.n32 VAPWR.n21 12.3338
R662 VAPWR.n28 VAPWR.n21 12.3338
R663 VAPWR.n8 VAPWR.n6 12.3338
R664 VAPWR.n11 VAPWR.n6 12.3338
R665 VAPWR.n9 VAPWR.n7 12.3338
R666 VAPWR.n12 VAPWR.n7 12.3338
R667 VAPWR.n78 VAPWR.n76 12.3338
R668 VAPWR.n92 VAPWR.n76 12.3338
R669 VAPWR.n77 VAPWR.n75 12.3338
R670 VAPWR.n91 VAPWR.n75 12.3338
R671 VAPWR.n66 VAPWR.n4 7.70883
R672 VAPWR.n60 VAPWR.n4 7.70883
R673 VAPWR.n118 VAPWR.n73 7.70883
R674 VAPWR.n112 VAPWR.n73 7.70883
R675 VAPWR.n125 VAPWR 4.11654
R676 VAPWR.n126 VAPWR 4.06671
R677 VAPWR.n123 VAPWR 3.16715
R678 VAPWR.n123 VAPWR 3.13288
R679 VAPWR.n39 VAPWR.n35 2.77496
R680 VAPWR.n39 VAPWR.n36 2.77496
R681 VAPWR.n50 VAPWR.n36 2.77496
R682 VAPWR.n22 VAPWR.n18 2.77496
R683 VAPWR.n22 VAPWR.n19 2.77496
R684 VAPWR.n33 VAPWR.n19 2.77496
R685 VAPWR.n16 VAPWR.n10 2.77496
R686 VAPWR.n17 VAPWR.n16 2.77496
R687 VAPWR.n98 VAPWR.n82 2.3255
R688 VAPWR.n108 VAPWR.n107 2.3255
R689 VAPWR.n54 VAPWR.n3 2.1216
R690 VAPWR.n89 VAPWR.n72 2.09672
R691 VAPWR.n52 VAPWR.n34 1.88425
R692 VAPWR.n106 VAPWR.n105 1.5505
R693 VAPWR.n10 VAPWR 1.40267
R694 VAPWR.n53 VAPWR.n52 1.37675
R695 VAPWR.n96 VAPWR.n95 1.32345
R696 VAPWR.n53 VAPWR.n17 1.23691
R697 VAPWR.n51 VAPWR.n50 1.22254
R698 VAPWR.n34 VAPWR.n33 1.22254
R699 VAPWR.n65 VAPWR.n1 1.163
R700 VAPWR.n117 VAPWR.n71 1.163
R701 VAPWR.n124 VAPWR.n123 1.07737
R702 VAPWR.n51 VAPWR.n35 0.894522
R703 VAPWR.n34 VAPWR.n18 0.894522
R704 VAPWR.n48 VAPWR.n35 0.845955
R705 VAPWR.n37 VAPWR.n36 0.845955
R706 VAPWR.n31 VAPWR.n18 0.845955
R707 VAPWR.n20 VAPWR.n19 0.845955
R708 VAPWR.n16 VAPWR.n15 0.845955
R709 VAPWR.n57 VAPWR.n56 0.845955
R710 VAPWR.n109 VAPWR.n108 0.845955
R711 VAPWR.t7 VAPWR.n63 0.81108
R712 VAPWR.t11 VAPWR.n115 0.81108
R713 VAPWR.n104 VAPWR.n103 0.797375
R714 VAPWR.n40 VAPWR.n39 0.664786
R715 VAPWR.n50 VAPWR.n49 0.664786
R716 VAPWR.n23 VAPWR.n22 0.664786
R717 VAPWR.n33 VAPWR.n32 0.664786
R718 VAPWR.n10 VAPWR.n9 0.664786
R719 VAPWR.n17 VAPWR.n8 0.664786
R720 VAPWR.n101 VAPWR.n78 0.664786
R721 VAPWR.n90 VAPWR.n77 0.664786
R722 VAPWR.n52 VAPWR.n51 0.5005
R723 VAPWR VAPWR.n126 0.491143
R724 VAPWR VAPWR.n88 0.490083
R725 VAPWR.n70 VAPWR.n1 0.448327
R726 VAPWR.n67 VAPWR.n66 0.404848
R727 VAPWR.n119 VAPWR.n118 0.404848
R728 VAPWR.n98 VAPWR.n97 0.3455
R729 VAPWR.n68 VAPWR.n0 0.313
R730 VAPWR.n125 VAPWR.n124 0.2968
R731 VAPWR.n103 VAPWR.n102 0.203625
R732 VAPWR.n96 VAPWR.n90 0.198256
R733 VAPWR.n70 VAPWR.n0 0.188
R734 VAPWR.n55 VAPWR.n54 0.179291
R735 VAPWR.n99 VAPWR.n98 0.163
R736 VAPWR.n56 VAPWR.n2 0.157262
R737 VAPWR.n119 VAPWR 0.152375
R738 VAPWR.n69 VAPWR.n68 0.143
R739 VAPWR.n101 VAPWR.n100 0.14175
R740 VAPWR.n70 VAPWR.n69 0.140949
R741 VAPWR VAPWR.n2 0.136533
R742 VAPWR.n104 VAPWR.n88 0.130708
R743 VAPWR VAPWR.n121 0.123855
R744 VAPWR VAPWR.n70 0.105837
R745 VAPWR.n90 VAPWR.n89 0.0951602
R746 VAPWR.n103 VAPWR.n101 0.0905
R747 VAPWR.n89 VAPWR.n79 0.0695895
R748 VAPWR.n121 VAPWR.n120 0.0690307
R749 VAPWR.n124 VAPWR 0.0651875
R750 VAPWR.n67 VAPWR.n2 0.062375
R751 VAPWR.n105 VAPWR 0.0568725
R752 VAPWR.n100 VAPWR.n99 0.0544216
R753 VAPWR.n122 VAPWR.n71 0.0533274
R754 VAPWR.n97 VAPWR 0.043
R755 VAPWR.n100 VAPWR 0.0364477
R756 VAPWR.n105 VAPWR 0.0364477
R757 VAPWR.n120 VAPWR.n119 0.033625
R758 VAPWR.n99 VAPWR.n96 0.0305
R759 VAPWR.n102 VAPWR 0.029875
R760 VAPWR.n56 VAPWR.n55 0.0297008
R761 VAPWR VAPWR.n122 0.0235263
R762 VAPWR VAPWR.n88 0.0212668
R763 VAPWR.n88 VAPWR 0.01927
R764 VAPWR VAPWR.n104 0.0184739
R765 VAPWR.n102 VAPWR 0.0152764
R766 VAPWR.n108 VAPWR.n79 0.0118818
R767 VAPWR.n108 VAPWR 0.00728914
R768 VAPWR.n122 VAPWR 0.00488596
R769 VAPWR.n54 VAPWR.n53 0.00425
R770 VAPWR.n126 VAPWR.n125 0.0033356
R771 VAPWR.n69 VAPWR.n67 0.002375
R772 flash_0.x2.clkb flash_0.x2.clkb.t0 167.038
R773 flash_0.x2.clkb flash_0.x2.clkb.t1 87.4292
R774 clk.n1 clk.t2 54.3383
R775 clk.n0 clk.t0 54.3383
R776 clk.n1 clk.t3 53.1307
R777 clk.n0 clk.t1 53.1307
R778 clk.n3 clk 39.2423
R779 clk.n3 clk.n2 9.04175
R780 clk.n2 clk 7.02925
R781 clk.n2 clk 3.72425
R782 clk clk.n1 0.2455
R783 clk clk.n0 0.2455
R784 clk clk.n3 0.078
R785 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t0 649.691
R786 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t1 227.442
R787 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t2 227.361
R788 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t5 216.731
R789 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t6 216.731
R790 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t3 216.731
R791 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t4 216.731
R792 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t7 216.731
R793 flash_0.x4.pos_mid_b flash_0.x4.pos_mid_b.t8 216.731
R794 ui_in[1].n0 ui_in[1].t17 207.43
R795 ui_in[1].n1 ui_in[1].t10 207.43
R796 ui_in[1].n2 ui_in[1].t12 207.43
R797 ui_in[1].n3 ui_in[1].t13 207.43
R798 ui_in[1].n4 ui_in[1].t15 207.43
R799 ui_in[1].n5 ui_in[1].t2 207.43
R800 ui_in[1].n26 ui_in[1].n23 123.867
R801 ui_in[1].n25 ui_in[1] 50.8126
R802 ui_in[1].n15 ui_in[1] 50.8126
R803 ui_in[1] ui_in[1].n1 48.5522
R804 ui_in[1] ui_in[1].n3 48.5522
R805 ui_in[1].n6 ui_in[1].n5 47.7953
R806 ui_in[1].n6 ui_in[1].n2 32.1435
R807 ui_in[1].n8 ui_in[1] 29.9794
R808 ui_in[1].n10 ui_in[1] 29.9794
R809 ui_in[1].n21 ui_in[1] 29.418
R810 ui_in[1].n18 ui_in[1] 29.418
R811 ui_in[1].n27 ui_in[1] 22.2876
R812 ui_in[1].n25 ui_in[1].n24 19.0005
R813 ui_in[1].n21 ui_in[1].n20 19.0005
R814 ui_in[1].n18 ui_in[1].n17 19.0005
R815 ui_in[1].n15 ui_in[1].n14 19.0005
R816 ui_in[1].n8 ui_in[1].n7 19.0005
R817 ui_in[1].n10 ui_in[1].n9 19.0005
R818 ui_in[1] ui_in[1].n0 13.6833
R819 ui_in[1] ui_in[1].n4 13.6833
R820 ui_in[1].n20 ui_in[1].t9 12.0505
R821 ui_in[1].n20 ui_in[1].t6 12.0505
R822 ui_in[1].n17 ui_in[1].t11 12.0505
R823 ui_in[1].n17 ui_in[1].t8 12.0505
R824 ui_in[1].n7 ui_in[1].t5 12.0505
R825 ui_in[1].n7 ui_in[1].t0 12.0505
R826 ui_in[1].n9 ui_in[1].t16 12.0505
R827 ui_in[1].n9 ui_in[1].t14 12.0505
R828 ui_in[1].n27 ui_in[1] 8.72144
R829 ui_in[1].n24 ui_in[1].t3 8.4355
R830 ui_in[1].n24 ui_in[1].t1 8.4355
R831 ui_in[1].n14 ui_in[1].t7 8.4355
R832 ui_in[1].n14 ui_in[1].t4 8.4355
R833 ui_in[1] ui_in[1].n26 4.94473
R834 ui_in[1].n13 ui_in[1].n12 4.5005
R835 ui_in[1].n2 ui_in[1] 3.75222
R836 ui_in[1].n1 ui_in[1] 3.75222
R837 ui_in[1].n0 ui_in[1] 3.75222
R838 ui_in[1].n5 ui_in[1] 3.75222
R839 ui_in[1].n4 ui_in[1] 3.75222
R840 ui_in[1].n3 ui_in[1] 3.75222
R841 ui_in[1].n28 ui_in[1].n13 3.61982
R842 ui_in[1].n11 ui_in[1].n8 2.96269
R843 ui_in[1].n12 ui_in[1].n6 1.69929
R844 ui_in[1].n16 ui_in[1].n15 1.59032
R845 ui_in[1].n22 ui_in[1].n19 1.42722
R846 ui_in[1].n19 ui_in[1].n18 1.32907
R847 ui_in[1].n22 ui_in[1].n21 1.32907
R848 ui_in[1].n26 ui_in[1].n25 1.32907
R849 ui_in[1].n11 ui_in[1].n10 1.32907
R850 ui_in[1].n23 ui_in[1].n16 1.29347
R851 ui_in[1].n12 ui_in[1].n11 0.48697
R852 ui_in[1].n19 ui_in[1].n16 0.25925
R853 ui_in[1].n23 ui_in[1].n22 0.25925
R854 ui_in[1].n13 ui_in[1] 0.0611061
R855 ui_in[1].n28 ui_in[1].n27 0.039875
R856 ui_in[1] ui_in[1].n28 0.0214375
R857 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t0 669.481
R858 flash_0.x4.neg_en_b.n0 flash_0.x4.neg_en_b.t1 669.481
R859 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t2 218.06
R860 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t3 218.06
R861 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t4 211.017
R862 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t6 208.394
R863 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t9 208.394
R864 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t5 207.43
R865 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t7 207.43
R866 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.t8 207.43
R867 flash_0.x4.neg_en_b flash_0.x4.neg_en_b.n0 50.3013
R868 flash_0.x4.neg_en_b.n0 flash_0.x4.neg_en_b 29.0914
R869 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t5 649.773
R870 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t4 649.691
R871 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.n1 594.383
R872 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.n2 594.301
R873 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t0 227.361
R874 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t8 216.731
R875 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t14 216.731
R876 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t13 216.731
R877 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.t9 105.956
R878 flash_0.x4.neg_mid_b.n0 flash_0.x4.neg_mid_b 103.529
R879 flash_0.x4.neg_mid_b.t8 flash_0.x4.neg_mid_b.t7 101.221
R880 flash_0.x4.neg_mid_b.t14 flash_0.x4.neg_mid_b.t12 101.221
R881 flash_0.x4.neg_mid_b.t13 flash_0.x4.neg_mid_b.t11 101.221
R882 flash_0.x4.neg_mid_b.n2 flash_0.x4.neg_mid_b.t3 55.3905
R883 flash_0.x4.neg_mid_b.n2 flash_0.x4.neg_mid_b.t6 55.3905
R884 flash_0.x4.neg_mid_b.n1 flash_0.x4.neg_mid_b.t1 55.3905
R885 flash_0.x4.neg_mid_b.n1 flash_0.x4.neg_mid_b.t2 55.3905
R886 flash_0.x4.neg_mid_b flash_0.x4.neg_mid_b.n0 23.6062
R887 flash_0.x4.neg_mid_b.n0 flash_0.x4.neg_mid_b.t10 22.3887
R888 flash_0.x4.dcgint.n0 flash_0.x4.dcgint.t8 644.461
R889 flash_0.x4.dcgint.n5 flash_0.x4.dcgint.t6 640.39
R890 flash_0.x4.dcgint.n3 flash_0.x4.dcgint.n1 605.365
R891 flash_0.x4.dcgint.n3 flash_0.x4.dcgint.n2 605.365
R892 flash_0.x4.dcgint.n4 flash_0.x4.dcgint.t5 477.228
R893 flash_0.x4.dcgint.t5 flash_0.x4.dcgint.t3 339.594
R894 flash_0.x4.dcgint.t3 flash_0.x4.dcgint.t9 339.594
R895 flash_0.x4.dcgint flash_0.x4.dcgint.t2 227.361
R896 flash_0.x4.dcgint flash_0.x4.dcgint.t1 227.361
R897 flash_0.x4.dcgint flash_0.x4.dcgint.t0 227.361
R898 flash_0.x4.dcgint.n4 flash_0.x4.dcgint.n3 69.5657
R899 flash_0.x4.dcgint.n1 flash_0.x4.dcgint.t4 55.3905
R900 flash_0.x4.dcgint.n1 flash_0.x4.dcgint.t10 55.3905
R901 flash_0.x4.dcgint.n2 flash_0.x4.dcgint.t7 55.3905
R902 flash_0.x4.dcgint.n2 flash_0.x4.dcgint.t11 55.3905
R903 flash_0.x4.dcgint.n6 flash_0.x4.dcgint.n5 9.3005
R904 flash_0.x4.dcgint.n5 flash_0.x4.dcgint.n4 8.9605
R905 flash_0.x4.dcgint flash_0.x4.dcgint.n6 7.52362
R906 flash_0.x4.dcgint.n6 flash_0.x4.dcgint.n0 1.14684
R907 flash_0.x4.dcgint.n4 flash_0.x4.dcgint.n0 1.0086
R908 flash_0.x7.pos_en_b.n1 flash_0.x7.pos_en_b.t0 669.481
R909 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b.t1 669.481
R910 flash_0.x7.pos_en_b flash_0.x7.pos_en_b.t2 218.06
R911 flash_0.x7.pos_en_b flash_0.x7.pos_en_b.t3 218.06
R912 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b.t6 65.4032
R913 flash_0.x7.pos_en_b.t6 flash_0.x7.pos_en_b 56.2429
R914 flash_0.x7.pos_en_b.t6 flash_0.x7.pos_en_b 56.2429
R915 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b 50.8126
R916 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b 50.8126
R917 flash_0.x7.pos_en_b flash_0.x7.pos_en_b.n1 29.0914
R918 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b 29.0914
R919 flash_0.x7.pos_en_b.n1 flash_0.x7.pos_en_b.n0 28.2591
R920 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b.t4 27.4355
R921 flash_0.x7.pos_en_b.n0 flash_0.x7.pos_en_b.t5 27.4355
R922 VDPWR.n84 VDPWR.n70 5586
R923 VDPWR.n84 VDPWR.n71 5586
R924 VDPWR.n79 VDPWR.n71 5586
R925 VDPWR.n79 VDPWR.n70 5586
R926 VDPWR.n129 VDPWR.n115 5586
R927 VDPWR.n129 VDPWR.n116 5586
R928 VDPWR.n124 VDPWR.n116 5586
R929 VDPWR.n124 VDPWR.n115 5586
R930 VDPWR.n30 VDPWR.n29 4689.72
R931 VDPWR.n27 VDPWR.n25 4689.72
R932 VDPWR.n80 VDPWR.n72 4509.29
R933 VDPWR.n125 VDPWR.n117 4509.29
R934 VDPWR.n83 VDPWR.n72 4506
R935 VDPWR.n128 VDPWR.n117 4506
R936 VDPWR.n44 VDPWR.n37 2442.35
R937 VDPWR.n41 VDPWR.n38 2442.35
R938 VDPWR.n61 VDPWR.n54 2442.35
R939 VDPWR.n58 VDPWR.n55 2442.35
R940 VDPWR.n83 VDPWR.t55 2271.78
R941 VDPWR.n128 VDPWR.t34 2271.78
R942 VDPWR.n30 VDPWR.n24 1828.1
R943 VDPWR.n28 VDPWR.n27 1828.1
R944 VDPWR.t22 VDPWR.t40 1429.17
R945 VDPWR.t38 VDPWR.t53 1429.17
R946 VDPWR.t55 VDPWR.n82 1226.56
R947 VDPWR.t34 VDPWR.n127 1226.56
R948 VDPWR.n26 VDPWR.n22 902.777
R949 VDPWR.n26 VDPWR.n23 902.777
R950 VDPWR.n31 VDPWR.n23 881.453
R951 VDPWR.n32 VDPWR.n22 879.466
R952 VDPWR.n33 VDPWR.t52 649.831
R953 VDPWR.n85 VDPWR.n69 627.201
R954 VDPWR.n78 VDPWR.n68 627.201
R955 VDPWR.n130 VDPWR.n114 627.201
R956 VDPWR.n123 VDPWR.n113 627.201
R957 VDPWR.n103 VDPWR.n102 585
R958 VDPWR.n98 VDPWR.n97 585
R959 VDPWR.n93 VDPWR.n92 585
R960 VDPWR.n101 VDPWR.n100 585
R961 VDPWR.n96 VDPWR.n95 585
R962 VDPWR.n91 VDPWR.n90 585
R963 VDPWR.n14 VDPWR.n13 585
R964 VDPWR.n9 VDPWR.n8 585
R965 VDPWR.n4 VDPWR.n3 585
R966 VDPWR.n12 VDPWR.n11 585
R967 VDPWR.n7 VDPWR.n6 585
R968 VDPWR.n2 VDPWR.n1 585
R969 VDPWR.n42 VDPWR.n37 535.419
R970 VDPWR.n43 VDPWR.n38 535.419
R971 VDPWR.n59 VDPWR.n54 535.419
R972 VDPWR.n60 VDPWR.n55 535.419
R973 VDPWR.n86 VDPWR.n85 525.553
R974 VDPWR.n131 VDPWR.n130 525.553
R975 VDPWR.n77 VDPWR.n69 492.048
R976 VDPWR.n122 VDPWR.n114 492.048
R977 VDPWR.n82 VDPWR.t22 394.779
R978 VDPWR.n127 VDPWR.t38 394.779
R979 VDPWR.n88 VDPWR.n66 297.151
R980 VDPWR.n107 VDPWR.n106 297.151
R981 VDPWR.n18 VDPWR.n17 297.151
R982 VDPWR.n111 VDPWR.n0 297.151
R983 VDPWR.n81 VDPWR.t30 272.363
R984 VDPWR.n126 VDPWR.t3 272.363
R985 VDPWR.n40 VDPWR.n36 260.519
R986 VDPWR.n45 VDPWR.n36 260.519
R987 VDPWR.n57 VDPWR.n53 260.519
R988 VDPWR.n62 VDPWR.n53 260.519
R989 VDPWR.n40 VDPWR.n39 232.66
R990 VDPWR.n46 VDPWR.n45 232.66
R991 VDPWR.n57 VDPWR.n56 232.66
R992 VDPWR.n63 VDPWR.n62 232.66
R993 VDPWR.n34 VDPWR.t12 228.215
R994 VDPWR.n51 VDPWR.t20 228.215
R995 VDPWR.t42 VDPWR.t32 172.133
R996 VDPWR.t36 VDPWR.t28 172.133
R997 VDPWR.t24 VDPWR.t36 172.133
R998 VDPWR.t30 VDPWR.t24 172.133
R999 VDPWR.t5 VDPWR.t9 172.133
R1000 VDPWR.t0 VDPWR.t13 172.133
R1001 VDPWR.t15 VDPWR.t0 172.133
R1002 VDPWR.t3 VDPWR.t15 172.133
R1003 VDPWR.n66 VDPWR.t23 160.44
R1004 VDPWR.n66 VDPWR.t56 160.44
R1005 VDPWR.n106 VDPWR.t27 160.44
R1006 VDPWR.n106 VDPWR.t41 160.44
R1007 VDPWR.n17 VDPWR.t8 160.44
R1008 VDPWR.n17 VDPWR.t54 160.44
R1009 VDPWR.n0 VDPWR.t39 160.44
R1010 VDPWR.n0 VDPWR.t35 160.44
R1011 VDPWR.n78 VDPWR.n77 135.154
R1012 VDPWR.n123 VDPWR.n122 135.154
R1013 VDPWR.t26 VDPWR.t42 135.093
R1014 VDPWR.t7 VDPWR.t5 135.093
R1015 VDPWR.n74 VDPWR 106.918
R1016 VDPWR.n119 VDPWR 106.918
R1017 VDPWR.n86 VDPWR.n68 101.647
R1018 VDPWR.n131 VDPWR.n113 101.647
R1019 VDPWR.n81 VDPWR.n80 57.7708
R1020 VDPWR.n126 VDPWR.n125 57.7708
R1021 VDPWR.n102 VDPWR.t25 55.3905
R1022 VDPWR.n102 VDPWR.t49 55.3905
R1023 VDPWR.n97 VDPWR.t47 55.3905
R1024 VDPWR.n97 VDPWR.t37 55.3905
R1025 VDPWR.n92 VDPWR.t33 55.3905
R1026 VDPWR.n92 VDPWR.t46 55.3905
R1027 VDPWR.n100 VDPWR.t48 55.3905
R1028 VDPWR.n100 VDPWR.t31 55.3905
R1029 VDPWR.n95 VDPWR.t29 55.3905
R1030 VDPWR.n95 VDPWR.t45 55.3905
R1031 VDPWR.n90 VDPWR.t50 55.3905
R1032 VDPWR.n90 VDPWR.t43 55.3905
R1033 VDPWR.n13 VDPWR.t57 55.3905
R1034 VDPWR.n13 VDPWR.t4 55.3905
R1035 VDPWR.n8 VDPWR.t14 55.3905
R1036 VDPWR.n8 VDPWR.t1 55.3905
R1037 VDPWR.n3 VDPWR.t17 55.3905
R1038 VDPWR.n3 VDPWR.t21 55.3905
R1039 VDPWR.n11 VDPWR.t16 55.3905
R1040 VDPWR.n11 VDPWR.t44 55.3905
R1041 VDPWR.n6 VDPWR.t18 55.3905
R1042 VDPWR.n6 VDPWR.t2 55.3905
R1043 VDPWR.n1 VDPWR.t10 55.3905
R1044 VDPWR.n1 VDPWR.t6 55.3905
R1045 VDPWR.t28 VDPWR.t26 37.0418
R1046 VDPWR.t13 VDPWR.t7 37.0418
R1047 VDPWR.n27 VDPWR.n26 37.0005
R1048 VDPWR.n31 VDPWR.n30 37.0005
R1049 VDPWR.n38 VDPWR.n36 30.8338
R1050 VDPWR.n37 VDPWR.n35 30.8338
R1051 VDPWR.n55 VDPWR.n53 30.8338
R1052 VDPWR.n54 VDPWR.n52 30.8338
R1053 VDPWR.n39 VDPWR.n35 27.8593
R1054 VDPWR.n46 VDPWR.n35 27.8593
R1055 VDPWR.n56 VDPWR.n52 27.8593
R1056 VDPWR.n63 VDPWR.n52 27.8593
R1057 VDPWR.n74 VDPWR.n73 19.0005
R1058 VDPWR.n119 VDPWR.n118 19.0005
R1059 VDPWR.n41 VDPWR.n40 16.8187
R1060 VDPWR.n45 VDPWR.n44 16.8187
R1061 VDPWR.n58 VDPWR.n57 16.8187
R1062 VDPWR.n62 VDPWR.n61 16.8187
R1063 VDPWR.n103 VDPWR 14.3064
R1064 VDPWR.n98 VDPWR 14.3064
R1065 VDPWR.n93 VDPWR 14.3064
R1066 VDPWR.n101 VDPWR 14.3064
R1067 VDPWR.n96 VDPWR 14.3064
R1068 VDPWR.n91 VDPWR 14.3064
R1069 VDPWR.n14 VDPWR 14.3064
R1070 VDPWR.n9 VDPWR 14.3064
R1071 VDPWR.n4 VDPWR 14.3064
R1072 VDPWR.n12 VDPWR 14.3064
R1073 VDPWR.n7 VDPWR 14.3064
R1074 VDPWR.n2 VDPWR 14.3064
R1075 VDPWR.n104 VDPWR.n103 13.8019
R1076 VDPWR.n99 VDPWR.n98 13.8019
R1077 VDPWR.n94 VDPWR.n93 13.8019
R1078 VDPWR.n104 VDPWR.n101 13.8019
R1079 VDPWR.n99 VDPWR.n96 13.8019
R1080 VDPWR.n94 VDPWR.n91 13.8019
R1081 VDPWR.n15 VDPWR.n14 13.8019
R1082 VDPWR.n10 VDPWR.n9 13.8019
R1083 VDPWR.n5 VDPWR.n4 13.8019
R1084 VDPWR.n15 VDPWR.n12 13.8019
R1085 VDPWR.n10 VDPWR.n7 13.8019
R1086 VDPWR.n5 VDPWR.n2 13.8019
R1087 VDPWR.n42 VDPWR.n41 13.0425
R1088 VDPWR.n44 VDPWR.n43 13.0425
R1089 VDPWR.n59 VDPWR.n58 13.0425
R1090 VDPWR.n61 VDPWR.n60 13.0425
R1091 VDPWR.t40 VDPWR.n81 10.895
R1092 VDPWR.t53 VDPWR.n126 10.895
R1093 VDPWR.n85 VDPWR.n84 10.2783
R1094 VDPWR.n84 VDPWR.n83 10.2783
R1095 VDPWR.n79 VDPWR.n78 10.2783
R1096 VDPWR.n80 VDPWR.n79 10.2783
R1097 VDPWR.n130 VDPWR.n129 10.2783
R1098 VDPWR.n129 VDPWR.n128 10.2783
R1099 VDPWR.n124 VDPWR.n123 10.2783
R1100 VDPWR.n125 VDPWR.n124 10.2783
R1101 VDPWR.n65 VDPWR.n64 9.74376
R1102 VDPWR.n39 VDPWR.n34 9.35589
R1103 VDPWR.n56 VDPWR.n51 9.35589
R1104 VDPWR VDPWR.n46 9.33194
R1105 VDPWR VDPWR.n63 9.33194
R1106 VDPWR.n73 VDPWR.t59 8.4355
R1107 VDPWR.n73 VDPWR.t58 8.4355
R1108 VDPWR.n118 VDPWR.t61 8.4355
R1109 VDPWR.n118 VDPWR.t60 8.4355
R1110 VDPWR.n70 VDPWR.n69 6.37981
R1111 VDPWR.n72 VDPWR.n70 6.37981
R1112 VDPWR.n71 VDPWR.n68 6.37981
R1113 VDPWR.n82 VDPWR.n71 6.37981
R1114 VDPWR.n115 VDPWR.n114 6.37981
R1115 VDPWR.n117 VDPWR.n115 6.37981
R1116 VDPWR.n116 VDPWR.n113 6.37981
R1117 VDPWR.n127 VDPWR.n116 6.37981
R1118 VDPWR.n48 VDPWR.n33 5.59737
R1119 VDPWR.n75 VDPWR.n67 4.51137
R1120 VDPWR.n120 VDPWR.n112 4.51137
R1121 VDPWR.n111 VDPWR.n110 3.96097
R1122 VDPWR.n89 VDPWR.n88 3.9605
R1123 VDPWR.n77 VDPWR.n76 3.88885
R1124 VDPWR.n122 VDPWR.n121 3.88885
R1125 VDPWR.n20 VDPWR 3.84311
R1126 VDPWR.n87 VDPWR.n67 3.7551
R1127 VDPWR.n132 VDPWR.n112 3.7551
R1128 VDPWR.n43 VDPWR.t11 3.68792
R1129 VDPWR.t11 VDPWR.n42 3.68792
R1130 VDPWR.n60 VDPWR.t19 3.68792
R1131 VDPWR.t19 VDPWR.n59 3.68792
R1132 VDPWR.n25 VDPWR.n22 3.03329
R1133 VDPWR.n29 VDPWR.n23 3.03329
R1134 VDPWR.n76 VDPWR.n74 2.3749
R1135 VDPWR.n121 VDPWR.n119 2.3749
R1136 VDPWR.n19 VDPWR.n18 2.25658
R1137 VDPWR.n108 VDPWR.n107 2.2555
R1138 VDPWR.n110 VDPWR.n19 1.98603
R1139 VDPWR.n33 VDPWR.n32 1.8605
R1140 VDPWR.n25 VDPWR.n24 1.85038
R1141 VDPWR.n29 VDPWR.n28 1.85038
R1142 VDPWR.n109 VDPWR.n108 1.7055
R1143 VDPWR.n49 VDPWR.n48 1.43592
R1144 VDPWR.n65 VDPWR.n50 1.29333
R1145 VDPWR.n28 VDPWR.t51 1.18321
R1146 VDPWR.t51 VDPWR.n24 1.18321
R1147 VDPWR.n32 VDPWR.n31 1.0245
R1148 VDPWR.n76 VDPWR.n75 0.813
R1149 VDPWR.n121 VDPWR.n120 0.813
R1150 VDPWR.n89 VDPWR.n65 0.683034
R1151 VDPWR.n85 VDPWR.n67 0.547559
R1152 VDPWR.n130 VDPWR.n112 0.547559
R1153 VDPWR.n48 VDPWR.n47 0.53175
R1154 VDPWR.n50 VDPWR.n49 0.486785
R1155 VDPWR.n110 VDPWR.n109 0.475641
R1156 VDPWR.n87 VDPWR.n86 0.4655
R1157 VDPWR.n132 VDPWR.n131 0.4655
R1158 VDPWR.n75 VDPWR.n69 0.344944
R1159 VDPWR.n120 VDPWR.n114 0.344944
R1160 VDPWR.n109 VDPWR.n89 0.278606
R1161 VDPWR.n19 VDPWR.n16 0.201021
R1162 VDPWR.n108 VDPWR.n105 0.182167
R1163 VDPWR.n21 VDPWR.n20 0.171
R1164 VDPWR.n107 VDPWR 0.102773
R1165 VDPWR.n18 VDPWR 0.102773
R1166 VDPWR.n99 VDPWR.n94 0.0902727
R1167 VDPWR.n10 VDPWR.n5 0.0902727
R1168 VDPWR.n105 VDPWR.n99 0.0772045
R1169 VDPWR.n16 VDPWR.n10 0.0772045
R1170 VDPWR.n21 VDPWR 0.0558125
R1171 VDPWR.n50 VDPWR.n20 0.0483835
R1172 VDPWR.n88 VDPWR 0.0483723
R1173 VDPWR VDPWR.n111 0.0483723
R1174 VDPWR.n47 VDPWR 0.0199611
R1175 VDPWR.n64 VDPWR 0.0199611
R1176 VDPWR.n49 VDPWR.n21 0.014875
R1177 VDPWR.n105 VDPWR.n104 0.0135682
R1178 VDPWR.n16 VDPWR.n15 0.0135682
R1179 VDPWR.n47 VDPWR.n34 0.00499102
R1180 VDPWR.n64 VDPWR.n51 0.00499102
R1181 VDPWR VDPWR.n87 0.00116489
R1182 VDPWR VDPWR.n132 0.00116489
R1183 ua[0].n6 ua[0].n4 2724.21
R1184 ua[0].n9 ua[0].n8 2724.21
R1185 ua[0].n7 ua[0].n6 1018.07
R1186 ua[0].n9 ua[0].n3 1018.07
R1187 ua[0].n12 ua[0].t3 649.886
R1188 ua[0].n0 ua[0].t1 649.692
R1189 ua[0].n5 ua[0].n1 526.307
R1190 ua[0].n5 ua[0].n2 526.307
R1191 ua[0].n10 ua[0].n2 497.486
R1192 ua[0].n11 ua[0].n1 493.762
R1193 ua[0].n6 ua[0].n5 37.0005
R1194 ua[0].n10 ua[0].n9 37.0005
R1195 ua[0].n14 ua[0] 13.435
R1196 ua[0].n4 ua[0].n1 5.78175
R1197 ua[0].n8 ua[0].n2 5.78175
R1198 ua[0].n0 ua[0].t0 4.69622
R1199 ua[0].n4 ua[0].n3 3.61407
R1200 ua[0].n8 ua[0].n7 3.61407
R1201 ua[0].t2 ua[0].n3 2.16152
R1202 ua[0].n7 ua[0].t2 2.16152
R1203 ua[0].n12 ua[0].n11 1.8605
R1204 ua[0].n11 ua[0].n10 1.54533
R1205 ua[0].n14 ua[0].n13 0.9005
R1206 ua[0].n13 ua[0].n0 0.64055
R1207 ua[0].n13 ua[0].n12 0.405262
R1208 ua[0] ua[0].n14 0.0639375
R1209 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t3 669.481
R1210 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t0 669.481
R1211 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t2 218.06
R1212 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t1 218.06
R1213 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t9 211.017
R1214 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t8 208.394
R1215 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t6 208.394
R1216 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t4 207.43
R1217 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t7 207.43
R1218 flash_0.x7.neg_en_b flash_0.x7.neg_en_b.t5 207.43
R1219 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t0 649.773
R1220 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t5 649.691
R1221 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.n3 594.383
R1222 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.n4 594.301
R1223 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t6 227.361
R1224 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t8 216.731
R1225 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t13 216.731
R1226 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.t14 216.731
R1227 flash_0.x7.neg_mid_b.n0 flash_0.x7.neg_mid_b.t15 105.956
R1228 flash_0.x7.neg_mid_b.n2 flash_0.x7.neg_mid_b 103.529
R1229 flash_0.x7.neg_mid_b.t8 flash_0.x7.neg_mid_b.t7 101.221
R1230 flash_0.x7.neg_mid_b.t13 flash_0.x7.neg_mid_b.t11 101.221
R1231 flash_0.x7.neg_mid_b.t14 flash_0.x7.neg_mid_b.t12 101.221
R1232 flash_0.x7.neg_mid_b.n4 flash_0.x7.neg_mid_b.t4 55.3905
R1233 flash_0.x7.neg_mid_b.n4 flash_0.x7.neg_mid_b.t2 55.3905
R1234 flash_0.x7.neg_mid_b.n3 flash_0.x7.neg_mid_b.t3 55.3905
R1235 flash_0.x7.neg_mid_b.n3 flash_0.x7.neg_mid_b.t1 55.3905
R1236 flash_0.x7.neg_mid_b.n2 flash_0.x7.neg_mid_b.n1 22.3887
R1237 flash_0.x7.neg_mid_b.n1 flash_0.x7.neg_mid_b.t10 8.4355
R1238 flash_0.x7.neg_mid_b.n1 flash_0.x7.neg_mid_b.t9 8.4355
R1239 flash_0.x7.neg_mid_b.n0 flash_0.x7.neg_mid_b 5.14452
R1240 flash_0.x7.neg_mid_b.n0 flash_0.x7.neg_mid_b.n2 2.45104
R1241 flash_0.x7.neg_mid_b flash_0.x7.neg_mid_b.n0 1.98963
R1242 flash_0.x6.Y flash_0.x6.Y.t0 228.901
R1243 flash_0.x5.A.n6 flash_0.x5.A.n4 2888.05
R1244 flash_0.x5.A.n9 flash_0.x5.A.n3 2888.05
R1245 flash_0.x5.A.n11 flash_0.x5.A.t3 658.039
R1246 flash_0.x5.A.n8 flash_0.x5.A.n4 509.978
R1247 flash_0.x5.A.n7 flash_0.x5.A.n3 509.978
R1248 flash_0.x5.A.n5 flash_0.x5.A.n2 334.683
R1249 flash_0.x5.A.n10 flash_0.x5.A.n2 334.683
R1250 flash_0.x5.A.n5 flash_0.x5.A.n1 291.084
R1251 flash_0.x5.A.n1 flash_0.x5.A.n10 290.635
R1252 flash_0.x5.A.n0 flash_0.x5.A.t0 215.056
R1253 flash_0.x5.A.n6 flash_0.x5.A.n5 146.25
R1254 flash_0.x5.A.n10 flash_0.x5.A.n9 146.25
R1255 flash_0.x5.A.n7 flash_0.x5.A.n6 114.621
R1256 flash_0.x5.A.n9 flash_0.x5.A.n8 114.621
R1257 flash_0.x5.A flash_0.x5.A.t4 33.6612
R1258 flash_0.x5.A flash_0.x5.A.t5 32.9049
R1259 flash_0.x5.A.n4 flash_0.x5.A.n2 32.5005
R1260 flash_0.x5.A.n3 flash_0.x5.A.n1 32.5005
R1261 flash_0.x5.A.t1 flash_0.x5.A.n7 25.8261
R1262 flash_0.x5.A.n8 flash_0.x5.A.t1 25.8261
R1263 flash_0.x5.A.n0 flash_0.x5.A.t2 17.2847
R1264 flash_0.x5.A flash_0.x5.A.n11 2.49814
R1265 flash_0.x5.A.n0 flash_0.x5.A.n1 1.43573
R1266 flash_0.x5.A.n11 flash_0.x5.A.n0 1.12981
R1267 ui_in[0].n0 ui_in[0].t6 207.43
R1268 ui_in[0].n1 ui_in[0].t14 207.43
R1269 ui_in[0].n2 ui_in[0].t8 207.43
R1270 ui_in[0].n3 ui_in[0].t9 207.43
R1271 ui_in[0].n4 ui_in[0].t0 207.43
R1272 ui_in[0].n5 ui_in[0].t10 207.43
R1273 ui_in[0].n26 ui_in[0].n23 123.867
R1274 ui_in[0].n25 ui_in[0] 50.8126
R1275 ui_in[0].n15 ui_in[0] 50.8126
R1276 ui_in[0] ui_in[0].n1 48.5522
R1277 ui_in[0] ui_in[0].n3 48.5522
R1278 ui_in[0].n6 ui_in[0].n5 47.7953
R1279 ui_in[0].n6 ui_in[0].n2 32.1435
R1280 ui_in[0].n8 ui_in[0] 29.9794
R1281 ui_in[0].n10 ui_in[0] 29.9794
R1282 ui_in[0].n21 ui_in[0] 29.418
R1283 ui_in[0].n18 ui_in[0] 29.418
R1284 ui_in[0].n27 ui_in[0] 26.7297
R1285 ui_in[0].n25 ui_in[0].n24 19.0005
R1286 ui_in[0].n21 ui_in[0].n20 19.0005
R1287 ui_in[0].n18 ui_in[0].n17 19.0005
R1288 ui_in[0].n15 ui_in[0].n14 19.0005
R1289 ui_in[0].n8 ui_in[0].n7 19.0005
R1290 ui_in[0].n10 ui_in[0].n9 19.0005
R1291 ui_in[0] ui_in[0].n0 13.6833
R1292 ui_in[0] ui_in[0].n4 13.6833
R1293 ui_in[0].n20 ui_in[0].t17 12.0505
R1294 ui_in[0].n20 ui_in[0].t15 12.0505
R1295 ui_in[0].n17 ui_in[0].t7 12.0505
R1296 ui_in[0].n17 ui_in[0].t4 12.0505
R1297 ui_in[0].n7 ui_in[0].t16 12.0505
R1298 ui_in[0].n7 ui_in[0].t12 12.0505
R1299 ui_in[0].n9 ui_in[0].t5 12.0505
R1300 ui_in[0].n9 ui_in[0].t2 12.0505
R1301 ui_in[0] ui_in[0].n13 11.4683
R1302 ui_in[0].n24 ui_in[0].t13 8.4355
R1303 ui_in[0].n24 ui_in[0].t11 8.4355
R1304 ui_in[0].n14 ui_in[0].t3 8.4355
R1305 ui_in[0].n14 ui_in[0].t1 8.4355
R1306 ui_in[0] ui_in[0].n26 4.94473
R1307 ui_in[0].n13 ui_in[0].n12 4.5005
R1308 ui_in[0].n13 ui_in[0] 4.0005
R1309 ui_in[0].n2 ui_in[0] 3.75222
R1310 ui_in[0].n1 ui_in[0] 3.75222
R1311 ui_in[0].n0 ui_in[0] 3.75222
R1312 ui_in[0].n5 ui_in[0] 3.75222
R1313 ui_in[0].n4 ui_in[0] 3.75222
R1314 ui_in[0].n3 ui_in[0] 3.75222
R1315 ui_in[0].n11 ui_in[0].n8 2.96269
R1316 ui_in[0].n27 ui_in[0] 2.12895
R1317 ui_in[0].n12 ui_in[0].n6 1.69929
R1318 ui_in[0].n16 ui_in[0].n15 1.59032
R1319 ui_in[0].n22 ui_in[0].n19 1.42722
R1320 ui_in[0].n19 ui_in[0].n18 1.32907
R1321 ui_in[0].n22 ui_in[0].n21 1.32907
R1322 ui_in[0].n26 ui_in[0].n25 1.32907
R1323 ui_in[0].n11 ui_in[0].n10 1.32907
R1324 ui_in[0].n23 ui_in[0].n16 1.29347
R1325 ui_in[0].n12 ui_in[0].n11 0.48697
R1326 ui_in[0].n19 ui_in[0].n16 0.25925
R1327 ui_in[0].n23 ui_in[0].n22 0.25925
R1328 ui_in[0].n13 ui_in[0] 0.0611061
R1329 ui_in[0] ui_in[0].n27 0.02925
R1330 flash_0.x7.VOUT.n8 flash_0.x7.VOUT.n6 2045.32
R1331 flash_0.x7.VOUT.n11 flash_0.x7.VOUT.n5 2045.32
R1332 flash_0.x7.VOUT.n9 flash_0.x7.VOUT.n8 836.909
R1333 flash_0.x7.VOUT.n11 flash_0.x7.VOUT.n10 836.909
R1334 flash_0.x7.VOUT flash_0.x7.VOUT.t4 649.691
R1335 flash_0.x7.VOUT flash_0.x7.VOUT.t10 649.691
R1336 flash_0.x7.VOUT flash_0.x7.VOUT.t11 649.691
R1337 flash_0.x7.VOUT flash_0.x7.VOUT.t6 649.691
R1338 flash_0.x7.VOUT flash_0.x7.VOUT.n2 594.383
R1339 flash_0.x7.VOUT flash_0.x7.VOUT.n13 594.301
R1340 flash_0.x7.VOUT flash_0.x7.VOUT.n14 594.301
R1341 flash_0.x7.VOUT flash_0.x7.VOUT.n3 594.301
R1342 flash_0.x7.VOUT flash_0.x7.VOUT.t7 227.431
R1343 flash_0.x7.VOUT flash_0.x7.VOUT.t8 227.361
R1344 flash_0.x7.VOUT.n6 flash_0.x7.VOUT.n4 195
R1345 flash_0.x7.VOUT.n12 flash_0.x7.VOUT.n11 146.25
R1346 flash_0.x7.VOUT.n8 flash_0.x7.VOUT.n7 146.25
R1347 flash_0.x7.VOUT.n12 flash_0.x7.VOUT.n4 132.894
R1348 flash_0.x7.VOUT.n7 flash_0.x7.VOUT.n4 132.894
R1349 flash_0.x7.VOUT.n9 flash_0.x7.VOUT.n5 105.183
R1350 flash_0.x7.VOUT.n10 flash_0.x7.VOUT.n6 105.183
R1351 flash_0.x7.VOUT.n12 flash_0.x7.VOUT.n1 53.1377
R1352 flash_0.x7.VOUT.n10 flash_0.x7.VOUT.t0 79.7913
R1353 flash_0.x7.VOUT.t0 flash_0.x7.VOUT.n9 79.7913
R1354 flash_0.x7.VOUT.n13 flash_0.x7.VOUT.t5 55.3905
R1355 flash_0.x7.VOUT.n13 flash_0.x7.VOUT.t3 55.3905
R1356 flash_0.x7.VOUT.n14 flash_0.x7.VOUT.t1 55.3905
R1357 flash_0.x7.VOUT.n14 flash_0.x7.VOUT.t2 55.3905
R1358 flash_0.x7.VOUT.n3 flash_0.x7.VOUT.t13 55.3905
R1359 flash_0.x7.VOUT.n3 flash_0.x7.VOUT.t12 55.3905
R1360 flash_0.x7.VOUT.n2 flash_0.x7.VOUT.t9 55.3905
R1361 flash_0.x7.VOUT.n2 flash_0.x7.VOUT.t14 55.3905
R1362 flash_0.x7.VOUT.n7 flash_0.x7.VOUT.n0 52.7987
R1363 flash_0.x7.VOUT flash_0.x7.VOUT.n0 28.5614
R1364 flash_0.x7.VOUT.n0 flash_0.x7.VOUT.n1 0.446827
R1365 flash_0.x7.VOUT.n5 flash_0.x7.VOUT.n1 198.951
R1366 w_7728_24730.t2 w_7728_24730.t0 336.07
R1367 w_7728_24730.t1 w_7728_24730.t2 649.856
R1368 w_7728_24730.t2 w_7728_24730.t3 649.692
R1369 flash_0.x3.clka flash_0.x3.clka.t0 167.038
R1370 flash_0.x3.clka flash_0.x3.clka.t1 87.4292
R1371 flash_0.x3.clkb flash_0.x3.clkb.t0 167.038
R1372 flash_0.x3.clkb flash_0.x3.clkb.t1 87.4292
R1373 flash_0.x4.pos_en_b.n0 flash_0.x4.pos_en_b.t0 669.481
R1374 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.t1 669.481
R1375 flash_0.x4.pos_en_b flash_0.x4.pos_en_b.t3 218.06
R1376 flash_0.x4.pos_en_b flash_0.x4.pos_en_b.t2 218.06
R1377 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.t4 65.4032
R1378 flash_0.x4.pos_en_b.t4 flash_0.x4.pos_en_b 56.2429
R1379 flash_0.x4.pos_en_b.t4 flash_0.x4.pos_en_b 56.2429
R1380 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b 50.8126
R1381 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b 50.8126
R1382 flash_0.x4.pos_en_b flash_0.x4.pos_en_b.n1 29.0914
R1383 flash_0.x4.pos_en_b.n0 flash_0.x4.pos_en_b 29.0914
R1384 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.n0 28.2591
R1385 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.t5 27.4355
R1386 flash_0.x4.pos_en_b.n1 flash_0.x4.pos_en_b.t6 27.4355
R1387 ui_in[2].n1 ui_in[2].t1 150.088
R1388 ui_in[2].n0 ui_in[2].t2 33.6007
R1389 ui_in[2].n0 ui_in[2].t0 32.9049
R1390 ui_in[2].n2 ui_in[2] 31.3871
R1391 ui_in[2].n2 ui_in[2].n1 4.55612
R1392 ui_in[2].n1 ui_in[2] 1.9712
R1393 ui_in[2] ui_in[2].n0 0.063
R1394 ui_in[2] ui_in[2].n2 0.047375
R1395 flash_0.x2.clka flash_0.x2.clka.t0 167.038
R1396 flash_0.x2.clka flash_0.x2.clka.t1 87.4292
R1397 flash_0.x7.dcgint.n0 flash_0.x7.dcgint.t4 644.461
R1398 flash_0.x7.dcgint.n5 flash_0.x7.dcgint.t1 640.39
R1399 flash_0.x7.dcgint.n3 flash_0.x7.dcgint.n1 605.365
R1400 flash_0.x7.dcgint.n3 flash_0.x7.dcgint.n2 605.365
R1401 flash_0.x7.dcgint.n4 flash_0.x7.dcgint.t0 477.228
R1402 flash_0.x7.dcgint.t0 flash_0.x7.dcgint.t2 339.594
R1403 flash_0.x7.dcgint.t2 flash_0.x7.dcgint.t6 339.594
R1404 flash_0.x7.dcgint flash_0.x7.dcgint.t11 227.361
R1405 flash_0.x7.dcgint flash_0.x7.dcgint.t10 227.361
R1406 flash_0.x7.dcgint flash_0.x7.dcgint.t9 227.361
R1407 flash_0.x7.dcgint.n4 flash_0.x7.dcgint.n3 69.5657
R1408 flash_0.x7.dcgint.n1 flash_0.x7.dcgint.t3 55.3905
R1409 flash_0.x7.dcgint.n1 flash_0.x7.dcgint.t7 55.3905
R1410 flash_0.x7.dcgint.n2 flash_0.x7.dcgint.t5 55.3905
R1411 flash_0.x7.dcgint.n2 flash_0.x7.dcgint.t8 55.3905
R1412 flash_0.x7.dcgint.n6 flash_0.x7.dcgint.n5 9.3005
R1413 flash_0.x7.dcgint.n5 flash_0.x7.dcgint.n4 8.9605
R1414 flash_0.x7.dcgint flash_0.x7.dcgint.n6 7.52362
R1415 flash_0.x7.dcgint.n6 flash_0.x7.dcgint.n0 1.14684
R1416 flash_0.x7.dcgint.n4 flash_0.x7.dcgint.n0 1.0086
R1417 uo_out[0].n0 uo_out[0].t0 228.901
R1418 uo_out[0].n0 uo_out[0].t1 84.4155
R1419 uo_out[0].n1 uo_out[0] 32.5825
R1420 uo_out[0].n1 uo_out[0].n0 4.88722
R1421 uo_out[0].n0 uo_out[0] 0.063
R1422 uo_out[0] uo_out[0].n1 0.016125
C0 flash_0.x4.neg_en_b flash_0.x4.neg_mid_b 0.430883f
C1 flash_0.x4.vintp flash_0.x4.pos_mid_b 0.252393f
C2 ui_in[0] flash_0.x4.VOUT 0.371415f
C3 flash_0.x5.A flash_0.x7.VPRGPOS 2.9732f
C4 flash_0.x4.neg_en_b ui_in[1] 3.07359f
C5 flash_0.x4.VOUT clk 0.069948f
C6 a_16296_28578# flash_0.x4.pos_en_b 3.62e-20
C7 flash_0.x7.dcgint ui_in[1] 0.239891f
C8 uo_out[0] flash_0.x7.VPRGNEG 3.06829f
C9 flash_0.x3.clkb flash_0.x3.clka 1.38778f
C10 flash_0.x4.VOUT flash_0.x7.VOUT 0.38054f
C11 flash_0.x4.VOUT flash_0.x2.clka 0.001465f
C12 flash_0.x4.pos_mid_b flash_0.x4.neg_mid_b 0.428431f
C13 ui_in[0] flash_0.x7.VDPWR1 0.001258f
C14 flash_0.x4.pos_mid flash_0.x4.neg_mid 4.98e-19
C15 ui_in[0] clk 4.50971f
C16 flash_0.x4.VOUT flash_0.x4.dcgint 0.619301f
C17 clk flash_0.x7.VDPWR1 2.14e-20
C18 flash_0.x3.clkb flash_0.x2.stage2 4.24817f
C19 flash_0.x4.neg_mid_b flash_0.x7.neg_mid_b 9.52e-20
C20 flash_0.x4.VOUT flash_0.x7.VPRGPOS 1.81837f
C21 flash_0.x4.pos_mid_b ui_in[1] 0.022428f
C22 uo_out[0] flash_0.x4.neg_en_b 0.00454f
C23 flash_0.x7.neg_mid a_20416_28577# 0.002271f
C24 ui_in[0] flash_0.x7.VOUT 0.473707f
C25 flash_0.x7.VDPWR1 flash_0.x7.VOUT 0.632531f
C26 flash_0.x4.pos_en_b flash_0.x4.neg_mid 0.080973f
C27 clk flash_0.x2.clka 0.357332f
C28 clk flash_0.x7.VOUT 2.11e-20
C29 uo_out[0] flash_0.x7.dcgint 0.003294f
C30 ui_in[1] flash_0.x7.neg_mid_b 0.208234f
C31 flash_0.x7.pos_mid_b flash_0.x4.neg_mid_b 4.26e-19
C32 flash_0.x7.neg_mid flash_0.x7.pos_en_b 0.080973f
C33 ui_in[0] flash_0.x4.dcgint 0.245012f
C34 ui_in[0] flash_0.x7.VPRGPOS 0.245007f
C35 flash_0.x2.clka flash_0.x7.VOUT 0.01934f
C36 flash_0.x4.pos_mid_b flash_0.x4.VDPWR1 0.264198f
C37 flash_0.x7.VDPWR1 flash_0.x7.VPRGPOS 1.29851f
C38 ui_in[1] flash_0.x7.pos_mid_b 0.773754f
C39 clk flash_0.x7.VPRGPOS 0.234475f
C40 flash_0.x7.VOUT flash_0.x4.dcgint 0.555359f
C41 flash_0.x2.clka flash_0.x7.VPRGPOS 0.589813f
C42 flash_0.x7.VOUT flash_0.x7.VPRGPOS 4.057f
C43 VDPWR a_7463_28281# 0.08485f
C44 flash_0.x2.clkinb flash_0.x2.stage1 0.189301f
C45 uo_out[0] flash_0.x7.neg_mid_b 0.030589f
C46 ui_in[2] a_7463_28281# 0.196624f
C47 VDPWR VAPWR 0.724319f
C48 VDPWR flash_0.x4.pos_mid 0.025715f
C49 flash_0.x4.dcgint flash_0.x7.VPRGPOS 0.026583f
C50 flash_0.x4.pos_mid ui_in[2] 0.022101f
C51 flash_0.x4.VOUT flash_0.x4.vintp 0.3705f
C52 VDPWR flash_0.x4.pos_en_b 1.86116f
C53 ui_in[2] flash_0.x4.pos_en_b 0.004173f
C54 ui_in[5] ui_in[6] 0.031023f
C55 flash_0.x4.VOUT flash_0.x4.neg_mid_b 0.500156f
C56 ui_in[0] flash_0.x4.vintp 8.2e-19
C57 ena clk 0.031023f
C58 VDPWR a_20416_28577# 0.106135f
C59 uo_out[0] flash_0.x5.A 0.225691f
C60 flash_0.x7.neg_mid_b flash_0.x7.pos_mid 3.38e-20
C61 flash_0.x4.VOUT ui_in[1] 0.456703f
C62 a_9352_28387# flash_0.x5.A 0.868312f
C63 VDPWR flash_0.x7.pos_en_b 1.80393f
C64 ui_in[0] flash_0.x4.neg_mid_b 0.209459f
C65 ui_in[2] flash_0.x7.pos_en_b 0.007039f
C66 clk flash_0.x4.neg_mid_b 2.05e-19
C67 flash_0.x4.vintp flash_0.x4.dcgint 1.54e-20
C68 flash_0.x7.pos_mid_b flash_0.x7.pos_mid 1.82667f
C69 flash_0.x4.vintp flash_0.x7.VPRGPOS 0.490137f
C70 flash_0.x4.VOUT flash_0.x4.VDPWR1 0.655265f
C71 ui_in[0] ui_in[1] 8.14454f
C72 flash_0.x7.VDPWR1 ui_in[1] 0.034551f
C73 ui_in[6] ui_in[7] 0.031023f
C74 flash_0.x7.VOUT flash_0.x4.neg_mid_b 0.002509f
C75 clk ui_in[1] 0.009319f
C76 flash_0.x3.clkb flash_0.x3.stage2 59.0307f
C77 VDPWR flash_0.x2.stage2 0.002548f
C78 flash_0.x4.VOUT uo_out[0] 0.031752f
C79 VDPWR flash_0.x2.clkb 0.024098f
C80 flash_0.x7.VPRGNEG VAPWR 2.20506f
C81 flash_0.x4.neg_mid_b flash_0.x4.dcgint 2.14914f
C82 flash_0.x4.VOUT a_9352_28387# 0.039663f
C83 ui_in[1] flash_0.x7.VOUT 0.636532f
C84 flash_0.x4.neg_mid_b flash_0.x7.VPRGPOS 0.008594f
C85 ui_in[0] flash_0.x4.VDPWR1 4.32e-20
C86 flash_0.x3.stage1 flash_0.x3.clkina 0.013783f
C87 clk flash_0.x4.VDPWR1 4.4e-19
C88 ui_in[1] flash_0.x4.dcgint 0.278517f
C89 flash_0.x4.VOUT flash_0.x2.stage1 3.9e-20
C90 flash_0.x3.stage1 flash_0.x3.clkinb 0.186066f
C91 flash_0.x7.VPRGNEG flash_0.x4.pos_en_b 0.232602f
C92 ui_in[0] uo_out[0] 0.016476f
C93 ui_in[1] flash_0.x7.VPRGPOS 0.63279f
C94 flash_0.x4.pos_mid flash_0.x4.neg_en_b 0.001081f
C95 uo_out[0] flash_0.x7.VOUT 0.093374f
C96 flash_0.x4.VDPWR1 flash_0.x4.dcgint 0.001075f
C97 flash_0.x7.VPRGNEG a_20416_28577# 0.062489f
C98 a_9352_28387# flash_0.x2.clka 0.002596f
C99 a_9352_28387# flash_0.x7.VOUT 0.834577f
C100 flash_0.x4.neg_en_b flash_0.x4.pos_en_b 0.337454f
C101 flash_0.x4.VDPWR1 flash_0.x7.VPRGPOS 1.31232f
C102 clk flash_0.x2.stage1 2.76362f
C103 flash_0.x2.clkinb VAPWR 1.65827f
C104 uo_out[0] flash_0.x4.dcgint 0.002825f
C105 flash_0.x7.VPRGNEG flash_0.x7.pos_en_b 0.22097f
C106 uo_out[0] flash_0.x7.VPRGPOS 2.61882f
C107 flash_0.x4.pos_mid flash_0.x4.pos_mid_b 1.82667f
C108 flash_0.x2.stage1 flash_0.x2.clka 57.610302f
C109 flash_0.x2.stage1 flash_0.x7.VOUT 0.001452f
C110 a_9352_28387# flash_0.x7.VPRGPOS 0.393793f
C111 flash_0.x4.vintp flash_0.x4.neg_mid_b 3.34e-19
C112 ui_in[0] flash_0.x7.pos_mid 7.01e-20
C113 uio_in[1] uio_in[2] 0.031023f
C114 clk flash_0.x7.pos_mid 8.13e-22
C115 flash_0.x4.neg_en_b flash_0.x7.pos_en_b 0.005326f
C116 flash_0.x7.VPRGNEG flash_0.x2.stage2 1.79888f
C117 flash_0.x4.pos_mid_b flash_0.x4.pos_en_b 0.391527f
C118 flash_0.x2.stage1 flash_0.x7.VPRGPOS 0.125764f
C119 flash_0.x2.clkb flash_0.x7.VPRGNEG 0.572269f
C120 flash_0.x7.neg_mid flash_0.x7.vintp 1.18e-20
C121 VAPWR flash_0.x3.clkina 1.05609f
C122 flash_0.x7.dcgint flash_0.x7.pos_en_b 0.178671f
C123 flash_0.x7.VOUT flash_0.x7.pos_mid 0.349932f
C124 VAPWR flash_0.x3.clkinb 1.66476f
C125 flash_0.x7.pos_mid flash_0.x4.dcgint 3.4e-19
C126 flash_0.x7.neg_mid flash_0.x7.neg_en_b 1.5384f
C127 ui_in[1] flash_0.x4.neg_mid_b 1.66762f
C128 flash_0.x4.vintp flash_0.x4.VDPWR1 0.235326f
C129 flash_0.x7.pos_mid flash_0.x7.VPRGPOS 0.417573f
C130 clk flash_0.x3.stage1 1.05122f
C131 a_20416_28577# flash_0.x7.neg_mid_b 0.166835f
C132 flash_0.x7.neg_mid_b flash_0.x7.pos_en_b 0.743046f
C133 flash_0.x2.clkinb flash_0.x2.stage2 0.359889f
C134 flash_0.x4.VDPWR1 flash_0.x4.neg_mid_b 0.00154f
C135 flash_0.x2.clkb flash_0.x2.clkinb 0.577668f
C136 uo_out[0] flash_0.x4.neg_mid_b 0.030267f
C137 flash_0.x7.pos_mid_b flash_0.x7.pos_en_b 0.391527f
C138 ui_in[1] flash_0.x4.VDPWR1 9.45e-21
C139 flash_0.x4.VOUT a_7463_28281# 0.069775f
C140 flash_0.x3.clka flash_0.x3.clkina 0.509107f
C141 flash_0.x3.clka flash_0.x3.clkinb 0.300643f
C142 uo_out[0] ui_in[1] 0.011391f
C143 flash_0.x4.VOUT flash_0.x4.pos_mid 0.012835f
C144 VDPWR flash_0.x7.vintp 0.003308f
C145 flash_0.x4.VOUT flash_0.x4.pos_en_b 0.142191f
C146 ui_in[2] flash_0.x7.vintp 0.007287f
C147 ui_in[0] flash_0.x4.pos_mid 0.343817f
C148 clk VAPWR 2.76692f
C149 flash_0.x4.pos_mid clk 1.68e-20
C150 flash_0.x4.neg_mid_b flash_0.x7.pos_mid 0.001667f
C151 flash_0.x2.clka a_7463_28281# 0.011214f
C152 a_7463_28281# flash_0.x7.VOUT 0.128388f
C153 VDPWR flash_0.x7.neg_en_b 1.678f
C154 ui_in[2] flash_0.x7.neg_en_b 0.010336f
C155 flash_0.x2.stage2 flash_0.x5.A 0.002905f
C156 flash_0.x2.clka VAPWR 0.417222f
C157 flash_0.x2.clkb flash_0.x5.A 0.05322f
C158 ui_in[0] flash_0.x4.pos_en_b 2.34221f
C159 ui_in[1] flash_0.x7.pos_mid 0.356278f
C160 clk flash_0.x4.pos_en_b 3.66e-19
C161 a_7463_28281# flash_0.x7.VPRGPOS 0.169831f
C162 a_16296_28578# flash_0.x4.neg_mid 0.002271f
C163 flash_0.x4.pos_mid flash_0.x7.VPRGPOS 0.416622f
C164 flash_0.x4.pos_en_b flash_0.x7.VOUT 0.023223f
C165 uio_in[3] uio_in[4] 0.031023f
C166 flash_0.x4.pos_en_b flash_0.x4.dcgint 0.178671f
C167 ui_in[0] flash_0.x7.pos_en_b 0.712549f
C168 flash_0.x7.VDPWR1 flash_0.x7.pos_en_b 4.17e-19
C169 flash_0.x4.pos_en_b flash_0.x7.VPRGPOS 0.064992f
C170 clk flash_0.x7.pos_en_b 1.99e-20
C171 a_20416_28577# flash_0.x7.VOUT 0.017698f
C172 clk flash_0.x3.clka 0.013936f
C173 flash_0.x7.VOUT flash_0.x7.pos_en_b 0.153015f
C174 flash_0.x7.pos_en_b flash_0.x4.dcgint 1.62e-19
C175 flash_0.x7.pos_en_b flash_0.x7.VPRGPOS 0.077604f
C176 flash_0.x2.stage2 flash_0.x2.clka 1.79536f
C177 flash_0.x4.pos_mid flash_0.x4.vintp 0.007513f
C178 flash_0.x2.stage2 flash_0.x7.VOUT 0.001251f
C179 flash_0.x7.VPRGNEG flash_0.x7.neg_en_b 0.007055f
C180 VDPWR a_16296_28578# 0.106132f
C181 flash_0.x2.clkb flash_0.x7.VOUT 0.084343f
C182 flash_0.x2.clkb flash_0.x2.clka 1.38778f
C183 flash_0.x2.clkinb flash_0.x2.clkina 0.886684f
C184 VDPWR ua[0] 0.053023f
C185 VDPWR flash_0.x7.neg_mid 1.38354f
C186 ui_in[2] ua[0] 0.009579f
C187 flash_0.x7.neg_mid ui_in[2] 0.001615f
C188 flash_0.x7.dcgint flash_0.x7.vintp 1.54e-20
C189 flash_0.x2.stage2 flash_0.x7.VPRGPOS 0.757314f
C190 flash_0.x4.vintp flash_0.x4.pos_en_b 0.014802f
C191 flash_0.x2.stage1 flash_0.x3.stage1 0.030249f
C192 flash_0.x2.clkb flash_0.x7.VPRGPOS 0.724895f
C193 flash_0.x3.stage2 flash_0.x3.clkina 0.20543f
C194 flash_0.x4.pos_mid flash_0.x4.neg_mid_b 3.38e-20
C195 flash_0.x3.stage2 flash_0.x3.clkinb 0.358189f
C196 flash_0.x7.dcgint flash_0.x7.neg_en_b 0.005849f
C197 VDPWR flash_0.x4.neg_mid 1.39258f
C198 flash_0.x4.pos_en_b flash_0.x4.neg_mid_b 0.743046f
C199 flash_0.x7.vintp flash_0.x7.neg_mid_b 3.34e-19
C200 ui_in[1] flash_0.x4.pos_en_b 0.711621f
C201 flash_0.x4.pos_mid flash_0.x4.VDPWR1 4.52e-20
C202 flash_0.x7.pos_mid_b flash_0.x7.vintp 0.252393f
C203 a_9352_28387# a_7463_28281# 0.06129f
C204 flash_0.x7.neg_mid_b flash_0.x7.neg_en_b 0.430883f
C205 flash_0.x4.neg_mid_b flash_0.x7.pos_en_b 1.35e-19
C206 ui_in[1] a_20416_28577# 2.08e-19
C207 flash_0.x4.VDPWR1 flash_0.x4.pos_en_b 4.58e-19
C208 VDPWR ua[7] 0.017072f
C209 flash_0.x7.VPRGNEG a_16296_28578# 0.062517f
C210 flash_0.x2.stage1 a_7463_28281# 1.01e-19
C211 flash_0.x7.pos_mid_b flash_0.x7.neg_en_b 0.013365f
C212 ui_in[1] flash_0.x7.pos_en_b 2.34386f
C213 uo_out[0] flash_0.x4.pos_en_b 0.012717f
C214 flash_0.x7.neg_mid flash_0.x7.VPRGNEG 0.976831f
C215 flash_0.x2.stage1 VAPWR 5.931509f
C216 ui_in[5] ui_in[4] 0.031023f
C217 flash_0.x2.stage2 flash_0.x4.neg_mid_b 0.002851f
C218 flash_0.x2.clkb flash_0.x4.neg_mid_b 7.35e-19
C219 VDPWR ui_in[2] 3.4924f
C220 flash_0.x4.neg_en_b a_16296_28578# 6.87e-21
C221 uo_out[0] a_20416_28577# 0.001639f
C222 flash_0.x7.VPRGNEG flash_0.x4.neg_mid 0.976831f
C223 flash_0.x7.neg_mid flash_0.x7.dcgint 1.61e-19
C224 uo_out[0] flash_0.x7.pos_en_b 0.01406f
C225 flash_0.x3.clkb flash_0.x3.clkina 0.005939f
C226 clk flash_0.x2.clkina 0.004029f
C227 uio_in[6] uio_in[7] 0.031023f
C228 flash_0.x3.clkb flash_0.x3.clkinb 0.57785f
C229 flash_0.x4.neg_en_b flash_0.x4.neg_mid 1.5384f
C230 uo_out[0] flash_0.x2.stage2 0.002424f
C231 flash_0.x3.stage2 flash_0.x7.VPRGPOS 1.93468f
C232 flash_0.x2.clka flash_0.x2.clkina 0.509107f
C233 uo_out[0] flash_0.x2.clkb 0.550211f
C234 flash_0.x2.stage1 flash_0.x3.clka 4.27357f
C235 flash_0.x3.stage1 VAPWR 4.90996f
C236 flash_0.x2.clkb a_9352_28387# 0.002716f
C237 ui_in[7] uio_in[0] 0.031023f
C238 flash_0.x7.VDPWR1 flash_0.x7.vintp 0.235326f
C239 flash_0.x7.neg_mid flash_0.x7.neg_mid_b 1.16207f
C240 flash_0.x7.VPRGPOS flash_0.x2.clkina 1.53e-19
C241 flash_0.x2.stage1 flash_0.x2.stage2 4.80565f
C242 flash_0.x2.clkb flash_0.x2.stage1 0.080777f
C243 flash_0.x7.pos_mid flash_0.x7.pos_en_b 0.595322f
C244 flash_0.x4.pos_mid_b flash_0.x4.neg_mid 0.001246f
C245 ui_in[0] flash_0.x7.neg_en_b 3.05692f
C246 flash_0.x7.neg_mid flash_0.x7.pos_mid_b 0.001246f
C247 flash_0.x7.VOUT flash_0.x7.vintp 0.396061f
C248 VDPWR flash_0.x7.VPRGNEG 13.5121f
C249 flash_0.x6.Y ua[0] 0.290173f
C250 flash_0.x7.VOUT flash_0.x7.neg_en_b 0.293369f
C251 flash_0.x7.vintp flash_0.x7.VPRGPOS 0.490248f
C252 VDPWR flash_0.x4.neg_en_b 1.82441f
C253 flash_0.x4.neg_en_b ui_in[2] 0.001238f
C254 VDPWR flash_0.x7.dcgint 0.006514f
C255 flash_0.x3.stage1 flash_0.x3.clka 57.6093f
C256 ui_in[2] flash_0.x7.dcgint 0.039612f
C257 ui_in[0] rst_n 0.031023f
C258 clk rst_n 0.031023f
C259 flash_0.x4.VOUT a_16296_28578# 0.017698f
C260 VDPWR flash_0.x4.pos_mid_b 0.038803f
C261 uio_in[3] uio_in[2] 0.031023f
C262 ui_in[2] flash_0.x4.pos_mid_b 0.047751f
C263 uio_in[1] uio_in[0] 0.031023f
C264 flash_0.x4.pos_mid flash_0.x4.pos_en_b 0.595322f
C265 VDPWR flash_0.x7.neg_mid_b 1.79805f
C266 ui_in[2] flash_0.x7.neg_mid_b 0.034018f
C267 ui_in[0] a_16296_28578# 2.08e-19
C268 flash_0.x3.clkb flash_0.x7.VPRGPOS 0.485638f
C269 VDPWR flash_0.x7.pos_mid_b 0.022461f
C270 ui_in[0] flash_0.x7.neg_mid 0.277486f
C271 flash_0.x4.VOUT flash_0.x4.neg_mid 0.069947f
C272 clk ua[0] 0.304224f
C273 ui_in[2] flash_0.x7.pos_mid_b 0.039178f
C274 VDPWR flash_0.x6.Y 7.946081f
C275 flash_0.x6.Y ui_in[2] 0.447688f
C276 uo_out[0] flash_0.x3.stage2 0.080392f
C277 flash_0.x7.neg_mid flash_0.x7.VOUT 0.070044f
C278 flash_0.x4.neg_en_b flash_0.x7.VPRGNEG 0.007732f
C279 VAPWR flash_0.x3.clka 1.5347f
C280 ui_in[1] flash_0.x7.vintp 0.004908f
C281 ui_in[0] flash_0.x4.neg_mid 0.003529f
C282 VDPWR flash_0.x5.A 2.1939f
C283 flash_0.x7.VPRGPOS ua[0] 0.043554f
C284 ui_in[2] flash_0.x5.A 0.032504f
C285 flash_0.x2.stage2 VAPWR 7.897181f
C286 flash_0.x7.neg_mid flash_0.x7.VPRGPOS 9.18e-20
C287 flash_0.x2.clkb VAPWR 0.392271f
C288 ui_in[1] flash_0.x7.neg_en_b 0.031249f
C289 flash_0.x7.VOUT flash_0.x4.neg_mid 1.16e-19
C290 flash_0.x2.stage1 flash_0.x2.clkina 0.01805f
C291 a_20416_28577# flash_0.x7.pos_en_b 3.62e-20
C292 flash_0.x7.VPRGNEG flash_0.x4.pos_mid_b 1.33e-19
C293 flash_0.x4.neg_mid flash_0.x4.dcgint 1.61e-19
C294 flash_0.x4.neg_mid flash_0.x7.VPRGPOS 1.81e-19
C295 uio_in[6] uio_in[5] 0.031023f
C296 flash_0.x7.VPRGNEG flash_0.x7.neg_mid_b 2.18563f
C297 flash_0.x4.VOUT VDPWR 1.92883f
C298 flash_0.x4.VOUT ui_in[2] 0.226315f
C299 uo_out[0] flash_0.x7.neg_en_b 0.00488f
C300 flash_0.x4.neg_en_b flash_0.x4.pos_mid_b 0.013365f
C301 flash_0.x7.VPRGNEG flash_0.x7.pos_mid_b 1.33e-19
C302 ui_in[0] VDPWR 3.54198f
C303 ui_in[3] ui_in[4] 0.031023f
C304 VDPWR flash_0.x7.VDPWR1 0.004126f
C305 ui_in[0] ui_in[2] 0.243794f
C306 VDPWR clk 0.460955f
C307 flash_0.x3.stage1 flash_0.x3.stage2 5.8896f
C308 flash_0.x7.VDPWR1 ui_in[2] 0.016435f
C309 clk ui_in[2] 2.12761f
C310 flash_0.x7.dcgint flash_0.x7.neg_mid_b 2.14914f
C311 flash_0.x2.stage2 flash_0.x3.clka 0.011129f
C312 uo_out[0] uio_in[7] 0.031023f
C313 flash_0.x7.vintp flash_0.x7.pos_mid 0.007513f
C314 a_16296_28578# flash_0.x4.neg_mid_b 0.166835f
C315 VDPWR flash_0.x7.VOUT 1.52997f
C316 ui_in[2] flash_0.x2.clka 0.003846f
C317 ui_in[2] flash_0.x7.VOUT 0.09898f
C318 flash_0.x2.clkb flash_0.x2.stage2 58.9902f
C319 flash_0.x7.dcgint flash_0.x7.pos_mid_b 0.009409f
C320 flash_0.x4.vintp flash_0.x4.neg_mid 1.18e-20
C321 VDPWR flash_0.x4.dcgint 0.046433f
C322 ui_in[2] flash_0.x4.dcgint 0.014403f
C323 flash_0.x7.pos_mid flash_0.x7.neg_en_b 0.001081f
C324 VDPWR flash_0.x7.VPRGPOS 1.07236f
C325 ui_in[2] flash_0.x7.VPRGPOS 0.388391f
C326 flash_0.x7.neg_mid ui_in[1] 0.003547f
C327 uio_in[5] uio_in[4] 0.031023f
C328 ui_in[3] ui_in[2] 0.031023f
C329 flash_0.x4.neg_mid_b flash_0.x4.neg_mid 1.16207f
C330 flash_0.x3.clkb flash_0.x2.stage1 7.28e-19
C331 flash_0.x4.VOUT flash_0.x7.VPRGNEG 0.387788f
C332 flash_0.x7.pos_mid_b flash_0.x7.neg_mid_b 0.428431f
C333 ui_in[1] flash_0.x4.neg_mid 0.277525f
C334 uo_out[0] a_16296_28578# 0.001641f
C335 VAPWR flash_0.x3.stage2 1.42027f
C336 flash_0.x7.neg_mid uo_out[0] 0.007637f
C337 flash_0.x3.clkinb flash_0.x3.clkina 0.886684f
C338 ui_in[0] flash_0.x7.VPRGNEG 0.063928f
C339 flash_0.x4.VOUT flash_0.x4.neg_en_b 0.293379f
C340 VDPWR flash_0.x4.vintp 0.003313f
C341 VAPWR flash_0.x2.clkina 1.04794f
C342 flash_0.x4.vintp ui_in[2] 0.00728f
C343 flash_0.x7.VPRGNEG flash_0.x7.VOUT 1.06096f
C344 uo_out[0] flash_0.x4.neg_mid 0.007647f
C345 ui_in[0] flash_0.x4.neg_en_b 0.030971f
C346 flash_0.x7.VPRGNEG flash_0.x4.dcgint 4.72e-19
C347 flash_0.x6.Y flash_0.x5.A 0.120397f
C348 ui_in[0] flash_0.x7.dcgint 0.146328f
C349 flash_0.x3.clkb flash_0.x3.stage1 0.07999f
C350 VDPWR flash_0.x4.neg_mid_b 1.91126f
C351 flash_0.x7.VDPWR1 flash_0.x7.dcgint 0.00211f
C352 flash_0.x4.VOUT flash_0.x4.pos_mid_b 0.255251f
C353 clk flash_0.x7.dcgint 2.23e-19
C354 flash_0.x7.VPRGNEG flash_0.x7.VPRGPOS 1.33754f
C355 ui_in[2] flash_0.x4.neg_mid_b 0.015154f
C356 flash_0.x4.neg_en_b flash_0.x7.VOUT 0.00256f
C357 flash_0.x7.neg_mid flash_0.x7.pos_mid 4.98e-19
C358 VDPWR ui_in[1] 3.6422f
C359 flash_0.x7.dcgint flash_0.x7.VOUT 0.61809f
C360 clk flash_0.x2.clkinb 0.350812f
C361 ui_in[2] ui_in[1] 4.33478f
C362 flash_0.x4.neg_en_b flash_0.x4.dcgint 0.005849f
C363 flash_0.x3.clka flash_0.x3.stage2 1.79536f
C364 ui_in[0] flash_0.x4.pos_mid_b 0.762651f
C365 flash_0.x4.neg_en_b flash_0.x7.VPRGPOS 0.002081f
C366 clk flash_0.x4.pos_mid_b 5.23e-19
C367 flash_0.x4.VOUT flash_0.x7.pos_mid_b 2.87e-22
C368 flash_0.x2.clkinb flash_0.x2.clka 0.30061f
C369 flash_0.x4.VOUT flash_0.x6.Y 0.044456f
C370 ui_in[0] flash_0.x7.neg_mid_b 1.58977f
C371 flash_0.x7.dcgint flash_0.x7.VPRGPOS 2.21e-19
C372 flash_0.x7.VDPWR1 flash_0.x7.neg_mid_b 0.0016f
C373 flash_0.x2.stage2 flash_0.x3.stage2 0.035345f
C374 VDPWR flash_0.x4.VDPWR1 0.004131f
C375 clk flash_0.x7.neg_mid_b 9.98e-21
C376 ui_in[2] flash_0.x4.VDPWR1 0.015856f
C377 flash_0.x4.pos_mid_b flash_0.x7.VOUT 5.14e-19
C378 VDPWR uo_out[0] 0.609895f
C379 flash_0.x2.clkinb flash_0.x7.VPRGPOS 2.41e-19
C380 ui_in[0] flash_0.x7.pos_mid_b 0.126143f
C381 flash_0.x4.pos_mid_b flash_0.x4.dcgint 0.009409f
C382 flash_0.x7.VDPWR1 flash_0.x7.pos_mid_b 0.264105f
C383 VDPWR a_9352_28387# 0.04147f
C384 flash_0.x7.VOUT flash_0.x7.neg_mid_b 0.501894f
C385 clk flash_0.x3.clkina 0.004029f
C386 uo_out[0] ui_in[2] 2.38891f
C387 clk flash_0.x7.pos_mid_b 2.14e-20
C388 flash_0.x2.stage2 flash_0.x2.clkina 0.206461f
C389 flash_0.x4.VOUT flash_0.x5.A 0.244704f
C390 flash_0.x2.clkb flash_0.x2.clkina 0.005816f
C391 flash_0.x4.pos_mid_b flash_0.x7.VPRGPOS 2.26733f
C392 flash_0.x7.vintp flash_0.x7.pos_en_b 0.014802f
C393 clk flash_0.x3.clkinb 0.350812f
C394 clk flash_0.x6.Y 0.154512f
C395 flash_0.x7.neg_mid_b flash_0.x4.dcgint 1.52e-19
C396 a_20416_28577# flash_0.x7.neg_en_b 6.87e-21
C397 flash_0.x7.pos_mid_b flash_0.x7.VOUT 0.781609f
C398 flash_0.x7.neg_mid_b flash_0.x7.VPRGPOS 0.003214f
C399 flash_0.x3.clkb VAPWR 0.370933f
C400 flash_0.x2.stage1 ui_in[2] 5.11e-19
C401 flash_0.x7.pos_en_b flash_0.x7.neg_en_b 0.337454f
C402 flash_0.x7.pos_mid_b flash_0.x4.dcgint 4.14e-19
C403 flash_0.x7.VPRGNEG flash_0.x4.neg_mid_b 2.19355f
C404 clk flash_0.x5.A 0.00419f
C405 flash_0.x7.pos_mid_b flash_0.x7.VPRGPOS 2.35676f
C406 flash_0.x6.Y flash_0.x7.VPRGPOS 0.054645f
C407 flash_0.x7.VPRGNEG ui_in[1] 0.065673f
C408 VDPWR flash_0.x7.pos_mid 0.018345f
C409 flash_0.x2.clka flash_0.x5.A 7.82e-19
C410 flash_0.x5.A flash_0.x7.VOUT 0.207778f
C411 ui_in[2] flash_0.x7.pos_mid 0.017392f
C412 ua[1] VGND 0.146962f
C413 ua[2] VGND 0.146962f
C414 ua[3] VGND 0.146962f
C415 ua[4] VGND 0.146962f
C416 ua[5] VGND 0.146962f
C417 ua[6] VGND 0.146962f
C418 ua[7] VGND 0.128006f
C419 ena VGND 0.070385f
C420 rst_n VGND 0.042875f
C421 ui_in[3] VGND 0.042875f
C422 ui_in[4] VGND 0.042875f
C423 ui_in[5] VGND 0.042875f
C424 ui_in[6] VGND 0.042875f
C425 ui_in[7] VGND 0.042875f
C426 uio_in[0] VGND 0.042875f
C427 uio_in[1] VGND 0.042875f
C428 uio_in[2] VGND 0.042875f
C429 uio_in[3] VGND 0.042875f
C430 uio_in[4] VGND 0.042875f
C431 uio_in[5] VGND 0.042875f
C432 uio_in[6] VGND 0.042875f
C433 uio_in[7] VGND 0.042875f
C434 ui_in[0] VGND 23.129925f
C435 ui_in[1] VGND 20.55118f
C436 uo_out[0] VGND 13.615086f
C437 ui_in[2] VGND 15.772717f
C438 clk VGND 25.498606f
C439 ua[0] VGND 35.369205f
C440 VDPWR VGND 96.2401f
C441 VAPWR VGND 43.180836f
C442 flash_0.x7.VDPWR1 VGND 0.460397f
C443 flash_0.x7.vintp VGND 0.039625f
C444 flash_0.x4.VDPWR1 VGND 0.472849f
C445 flash_0.x4.vintp VGND 0.051188f
C446 flash_0.x7.pos_mid VGND 1.29059f
C447 flash_0.x7.pos_mid_b VGND 3.896975f
C448 flash_0.x4.pos_mid VGND 1.31994f
C449 flash_0.x4.pos_mid_b VGND 3.985879f
C450 flash_0.x6.Y VGND 13.697189f
C451 flash_0.x7.neg_en_b VGND 3.319393f
C452 flash_0.x7.neg_mid VGND 0.210934f
C453 a_20416_28577# VGND 0.048706f
C454 flash_0.x7.neg_mid_b VGND 4.319581f
C455 flash_0.x7.pos_en_b VGND 7.747194f
C456 flash_0.x4.neg_en_b VGND 3.199902f
C457 flash_0.x4.neg_mid VGND 0.206959f
C458 a_16296_28578# VGND 0.047639f
C459 flash_0.x4.neg_mid_b VGND 4.854208f
C460 flash_0.x4.pos_en_b VGND 7.770404f
C461 a_9352_28387# VGND 0.21567f
C462 flash_0.x4.VOUT VGND 4.498701f
C463 a_7463_28281# VGND 0.801294f
C464 flash_0.x2.clkb VGND 63.13064f
C465 flash_0.x2.clka VGND 62.52466f
C466 flash_0.x2.clkinb VGND 3.11026f
C467 flash_0.x2.clkina VGND 1.57797f
C468 flash_0.x3.clkb VGND 66.16767f
C469 flash_0.x3.clka VGND 65.171394f
C470 flash_0.x3.clkinb VGND 3.10612f
C471 flash_0.x3.clkina VGND 1.5755f
C472 flash_0.x7.dcgint VGND 3.309877f
C473 flash_0.x4.dcgint VGND 2.988657f
C474 flash_0.x5.A VGND 5.742692f
C475 flash_0.x7.VOUT VGND 11.406838f
C476 flash_0.x7.VPRGNEG VGND 80.182205f
C477 flash_0.x2.stage2 VGND 15.4695f
C478 flash_0.x2.stage1 VGND 18.413f
C479 flash_0.x7.VPRGPOS VGND 0.145575p
C480 flash_0.x3.stage2 VGND 24.3058f
C481 flash_0.x3.stage1 VGND 23.173801f
C482 uo_out[0].t0 VGND 0.038292f
C483 uo_out[0].t1 VGND 0.037022f
C484 uo_out[0].n0 VGND 0.257992f
C485 uo_out[0].n1 VGND 3.39873f
C486 flash_0.x7.dcgint.t9 VGND 0.016015f
C487 flash_0.x7.dcgint.t10 VGND 0.016015f
C488 flash_0.x7.dcgint.t11 VGND 0.016015f
C489 flash_0.x7.dcgint.t4 VGND 0.017561f
C490 flash_0.x7.dcgint.n0 VGND 0.05401f
C491 flash_0.x7.dcgint.t1 VGND 0.017266f
C492 flash_0.x7.dcgint.t6 VGND 0.355987f
C493 flash_0.x7.dcgint.t2 VGND 0.222316f
C494 flash_0.x7.dcgint.t0 VGND 0.280884f
C495 flash_0.x7.dcgint.t3 VGND 0.004616f
C496 flash_0.x7.dcgint.t7 VGND 0.004616f
C497 flash_0.x7.dcgint.n1 VGND 0.009325f
C498 flash_0.x7.dcgint.t5 VGND 0.004616f
C499 flash_0.x7.dcgint.t8 VGND 0.004616f
C500 flash_0.x7.dcgint.n2 VGND 0.009325f
C501 flash_0.x7.dcgint.n3 VGND 0.045712f
C502 flash_0.x7.dcgint.n4 VGND 0.233815f
C503 flash_0.x7.dcgint.n5 VGND 0.046322f
C504 flash_0.x7.dcgint.n6 VGND 0.34091f
C505 flash_0.x2.clka.t1 VGND 0.011299f
C506 flash_0.x2.clka.t0 VGND 0.017732f
C507 ui_in[2].t2 VGND 0.727097f
C508 ui_in[2].t0 VGND 0.69579f
C509 ui_in[2].n0 VGND 0.550323f
C510 ui_in[2].t1 VGND 0.186184f
C511 ui_in[2].n1 VGND 1.11593f
C512 ui_in[2].n2 VGND 4.46526f
C513 flash_0.x4.pos_en_b.n0 VGND 0.032452f
C514 flash_0.x4.pos_en_b.n1 VGND 0.766491f
C515 flash_0.x4.pos_en_b.t4 VGND 0.932199f
C516 flash_0.x4.pos_en_b.t5 VGND 0.216253f
C517 flash_0.x4.pos_en_b.t6 VGND 0.216253f
C518 flash_0.x4.pos_en_b.t1 VGND 0.010089f
C519 flash_0.x4.pos_en_b.t0 VGND 0.010089f
C520 flash_0.x4.pos_en_b.t2 VGND 0.008975f
C521 flash_0.x4.pos_en_b.t3 VGND 0.008975f
C522 flash_0.x3.clkb.t1 VGND 0.012451f
C523 flash_0.x3.clkb.t0 VGND 0.01954f
C524 flash_0.x3.clka.t1 VGND 0.012142f
C525 flash_0.x3.clka.t0 VGND 0.019055f
C526 w_7728_24730.t0 VGND 6.5007f
C527 w_7728_24730.t2 VGND 6.37557f
C528 w_7728_24730.t3 VGND 0.011863f
C529 w_7728_24730.t1 VGND 0.01187f
C530 flash_0.x7.VOUT.n0 VGND 1.34521f
C531 flash_0.x7.VOUT.n1 VGND 0.023832f
C532 flash_0.x7.VOUT.t11 VGND 0.009996f
C533 flash_0.x7.VOUT.t9 VGND 0.002635f
C534 flash_0.x7.VOUT.t14 VGND 0.002635f
C535 flash_0.x7.VOUT.n2 VGND 0.005414f
C536 flash_0.x7.VOUT.t13 VGND 0.002635f
C537 flash_0.x7.VOUT.t12 VGND 0.002635f
C538 flash_0.x7.VOUT.n3 VGND 0.005412f
C539 flash_0.x7.VOUT.t10 VGND 0.009996f
C540 flash_0.x7.VOUT.t7 VGND 0.009046f
C541 flash_0.x7.VOUT.t8 VGND 0.009042f
C542 flash_0.x7.VOUT.n4 VGND 0.02291f
C543 flash_0.x7.VOUT.n5 VGND 0.02319f
C544 flash_0.x7.VOUT.n6 VGND 0.02291f
C545 flash_0.x7.VOUT.n7 VGND 0.017131f
C546 flash_0.x7.VOUT.n8 VGND 0.148335f
C547 flash_0.x7.VOUT.t0 VGND 0.1867f
C548 flash_0.x7.VOUT.n11 VGND 0.148335f
C549 flash_0.x7.VOUT.n12 VGND 0.016888f
C550 flash_0.x7.VOUT.t6 VGND 0.009331f
C551 flash_0.x7.VOUT.t4 VGND 0.009331f
C552 flash_0.x7.VOUT.t5 VGND 0.002635f
C553 flash_0.x7.VOUT.t3 VGND 0.002635f
C554 flash_0.x7.VOUT.n13 VGND 0.005412f
C555 flash_0.x7.VOUT.t1 VGND 0.002635f
C556 flash_0.x7.VOUT.t2 VGND 0.002635f
C557 flash_0.x7.VOUT.n14 VGND 0.005412f
C558 ui_in[0].t6 VGND 0.037781f
C559 ui_in[0].n0 VGND 0.057717f
C560 ui_in[0].t14 VGND 0.037781f
C561 ui_in[0].n1 VGND 0.14905f
C562 ui_in[0].t8 VGND 0.037781f
C563 ui_in[0].n2 VGND 0.109725f
C564 ui_in[0].t9 VGND 0.037781f
C565 ui_in[0].n3 VGND 0.14905f
C566 ui_in[0].t0 VGND 0.037781f
C567 ui_in[0].n4 VGND 0.057717f
C568 ui_in[0].t10 VGND 0.037781f
C569 ui_in[0].n5 VGND 0.146838f
C570 ui_in[0].n6 VGND 0.408027f
C571 ui_in[0].t16 VGND 0.266104f
C572 ui_in[0].t12 VGND 0.278064f
C573 ui_in[0].n7 VGND 0.44849f
C574 ui_in[0].n8 VGND 0.330488f
C575 ui_in[0].t5 VGND 0.266104f
C576 ui_in[0].t2 VGND 0.278064f
C577 ui_in[0].n9 VGND 0.44849f
C578 ui_in[0].n10 VGND 0.227519f
C579 ui_in[0].n11 VGND 0.226122f
C580 ui_in[0].n12 VGND 0.127227f
C581 ui_in[0].n13 VGND 1.01912f
C582 ui_in[0].t3 VGND 0.22275f
C583 ui_in[0].t1 VGND 0.20481f
C584 ui_in[0].n14 VGND 0.313943f
C585 ui_in[0].n15 VGND 0.120049f
C586 ui_in[0].n16 VGND 0.1624f
C587 ui_in[0].t7 VGND 0.266104f
C588 ui_in[0].t4 VGND 0.278064f
C589 ui_in[0].n17 VGND 0.44849f
C590 ui_in[0].n18 VGND 0.223258f
C591 ui_in[0].n19 VGND 0.099266f
C592 ui_in[0].t17 VGND 0.266104f
C593 ui_in[0].t15 VGND 0.278064f
C594 ui_in[0].n20 VGND 0.44849f
C595 ui_in[0].n21 VGND 0.223258f
C596 ui_in[0].n22 VGND 0.099844f
C597 ui_in[0].n23 VGND 0.313671f
C598 ui_in[0].t13 VGND 0.22275f
C599 ui_in[0].t11 VGND 0.20481f
C600 ui_in[0].n24 VGND 0.313943f
C601 ui_in[0].n25 VGND 0.129255f
C602 ui_in[0].n26 VGND 0.508238f
C603 ui_in[0].n27 VGND 3.80721f
C604 flash_0.x5.A.n0 VGND 0.493086f
C605 flash_0.x5.A.n1 VGND 0.103919f
C606 flash_0.x5.A.t5 VGND 0.417187f
C607 flash_0.x5.A.t4 VGND 0.436255f
C608 flash_0.x5.A.t3 VGND 0.014943f
C609 flash_0.x5.A.n2 VGND 0.065317f
C610 flash_0.x5.A.n3 VGND 0.639596f
C611 flash_0.x5.A.n4 VGND 0.639596f
C612 flash_0.x5.A.n5 VGND 0.068344f
C613 flash_0.x5.A.n6 VGND 0.114375f
C614 flash_0.x5.A.t1 VGND 0.747064f
C615 flash_0.x5.A.n9 VGND 0.114375f
C616 flash_0.x5.A.n10 VGND 0.06833f
C617 flash_0.x5.A.t2 VGND 0.110389f
C618 flash_0.x5.A.t0 VGND 0.169707f
C619 flash_0.x5.A.n11 VGND 0.595547f
C620 flash_0.x6.Y.t0 VGND 0.039316f
C621 flash_0.x7.neg_mid_b.n0 VGND 0.539196f
C622 flash_0.x7.neg_mid_b.t10 VGND 0.243062f
C623 flash_0.x7.neg_mid_b.t9 VGND 0.243062f
C624 flash_0.x7.neg_mid_b.n1 VGND 0.341911f
C625 flash_0.x7.neg_mid_b.n2 VGND 0.140489f
C626 flash_0.x7.neg_mid_b.t0 VGND 0.027096f
C627 flash_0.x7.neg_mid_b.t3 VGND 0.007678f
C628 flash_0.x7.neg_mid_b.t1 VGND 0.007678f
C629 flash_0.x7.neg_mid_b.n3 VGND 0.015666f
C630 flash_0.x7.neg_mid_b.t15 VGND 0.085863f
C631 flash_0.x7.neg_mid_b.t6 VGND 0.02816f
C632 flash_0.x7.neg_mid_b.t7 VGND 0.067252f
C633 flash_0.x7.neg_mid_b.t8 VGND 0.122491f
C634 flash_0.x7.neg_mid_b.t11 VGND 0.067252f
C635 flash_0.x7.neg_mid_b.t13 VGND 0.122491f
C636 flash_0.x7.neg_mid_b.t12 VGND 0.067252f
C637 flash_0.x7.neg_mid_b.t14 VGND 0.122491f
C638 flash_0.x7.neg_mid_b.t4 VGND 0.007678f
C639 flash_0.x7.neg_mid_b.t2 VGND 0.007678f
C640 flash_0.x7.neg_mid_b.n4 VGND 0.015661f
C641 flash_0.x7.neg_mid_b.t5 VGND 0.02709f
C642 flash_0.x7.neg_en_b.t0 VGND 0.038945f
C643 flash_0.x7.neg_en_b.t9 VGND 0.052338f
C644 flash_0.x7.neg_en_b.t5 VGND 0.051225f
C645 flash_0.x7.neg_en_b.t7 VGND 0.051225f
C646 flash_0.x7.neg_en_b.t4 VGND 0.051225f
C647 flash_0.x7.neg_en_b.t8 VGND 0.051201f
C648 flash_0.x7.neg_en_b.t6 VGND 0.051201f
C649 flash_0.x7.neg_en_b.t3 VGND 0.036466f
C650 flash_0.x7.neg_en_b.t1 VGND 0.032439f
C651 flash_0.x7.neg_en_b.t2 VGND 0.032439f
C652 ua[0].t1 VGND 0.00285f
C653 ua[0].t0 VGND 0.716764f
C654 ua[0].n0 VGND 0.259475f
C655 ua[0].t3 VGND 0.002851f
C656 ua[0].n1 VGND 0.024193f
C657 ua[0].n2 VGND 0.02427f
C658 ua[0].n4 VGND 0.042071f
C659 ua[0].n5 VGND 0.02521f
C660 ua[0].n6 VGND 0.281781f
C661 ua[0].t2 VGND 0.430674f
C662 ua[0].n8 VGND 0.042071f
C663 ua[0].n9 VGND 0.281781f
C664 ua[0].n10 VGND 0.015559f
C665 ua[0].n11 VGND 0.0156f
C666 ua[0].n12 VGND -0.00395f
C667 ua[0].n13 VGND 0.015585f
C668 ua[0].n14 VGND 1.92631f
C669 VDPWR.t39 VGND 0.003648f
C670 VDPWR.t35 VGND 0.003648f
C671 VDPWR.n0 VGND 0.007478f
C672 VDPWR.t10 VGND 0.001259f
C673 VDPWR.t6 VGND 0.001259f
C674 VDPWR.n1 VGND 0.002519f
C675 VDPWR.n2 VGND 0.003602f
C676 VDPWR.t17 VGND 0.001259f
C677 VDPWR.t21 VGND 0.001259f
C678 VDPWR.n3 VGND 0.002519f
C679 VDPWR.n4 VGND 0.003602f
C680 VDPWR.n5 VGND 0.076297f
C681 VDPWR.t18 VGND 0.001259f
C682 VDPWR.t2 VGND 0.001259f
C683 VDPWR.n6 VGND 0.002519f
C684 VDPWR.n7 VGND 0.003602f
C685 VDPWR.t14 VGND 0.001259f
C686 VDPWR.t1 VGND 0.001259f
C687 VDPWR.n8 VGND 0.002519f
C688 VDPWR.n9 VGND 0.003602f
C689 VDPWR.n10 VGND 0.117955f
C690 VDPWR.t16 VGND 0.001259f
C691 VDPWR.t44 VGND 0.001259f
C692 VDPWR.n11 VGND 0.002519f
C693 VDPWR.n12 VGND 0.003602f
C694 VDPWR.t57 VGND 0.001259f
C695 VDPWR.t4 VGND 0.001259f
C696 VDPWR.n13 VGND 0.002519f
C697 VDPWR.n14 VGND 0.003602f
C698 VDPWR.n15 VGND 0.024702f
C699 VDPWR.n16 VGND 0.074832f
C700 VDPWR.t8 VGND 0.003648f
C701 VDPWR.t54 VGND 0.003648f
C702 VDPWR.n17 VGND 0.007478f
C703 VDPWR.n18 VGND 0.020625f
C704 VDPWR.n19 VGND 0.047136f
C705 VDPWR.n20 VGND 10.0402f
C706 VDPWR.n21 VGND 0.037822f
C707 VDPWR.t52 VGND 0.004764f
C708 VDPWR.n22 VGND 0.070102f
C709 VDPWR.n23 VGND 0.070176f
C710 VDPWR.n25 VGND 0.120477f
C711 VDPWR.n26 VGND 0.071725f
C712 VDPWR.n27 VGND 0.823306f
C713 VDPWR.t51 VGND 1.32138f
C714 VDPWR.n29 VGND 0.120477f
C715 VDPWR.n30 VGND 0.823306f
C716 VDPWR.n31 VGND 0.03915f
C717 VDPWR.n32 VGND 0.039161f
C718 VDPWR.n33 VGND 0.298525f
C719 VDPWR.t12 VGND 0.009255f
C720 VDPWR.n34 VGND 0.02185f
C721 VDPWR.n35 VGND 0.002185f
C722 VDPWR.n36 VGND 0.021079f
C723 VDPWR.n37 VGND 0.166406f
C724 VDPWR.n38 VGND 0.166406f
C725 VDPWR.n39 VGND 0.010632f
C726 VDPWR.n40 VGND 0.019667f
C727 VDPWR.n41 VGND 0.020798f
C728 VDPWR.t11 VGND 0.259082f
C729 VDPWR.n44 VGND 0.020798f
C730 VDPWR.n45 VGND 0.019667f
C731 VDPWR.n46 VGND 0.010601f
C732 VDPWR.n47 VGND 0.031206f
C733 VDPWR.n48 VGND 0.366962f
C734 VDPWR.n49 VGND 0.117793f
C735 VDPWR.n50 VGND 0.840951f
C736 VDPWR.t20 VGND 0.009255f
C737 VDPWR.n51 VGND 0.02185f
C738 VDPWR.n52 VGND 0.002185f
C739 VDPWR.n53 VGND 0.021079f
C740 VDPWR.n54 VGND 0.166406f
C741 VDPWR.n55 VGND 0.166406f
C742 VDPWR.n56 VGND 0.010632f
C743 VDPWR.n57 VGND 0.019667f
C744 VDPWR.n58 VGND 0.020798f
C745 VDPWR.t19 VGND 0.259082f
C746 VDPWR.n61 VGND 0.020798f
C747 VDPWR.n62 VGND 0.019667f
C748 VDPWR.n63 VGND 0.010601f
C749 VDPWR.n64 VGND 0.076647f
C750 VDPWR.n65 VGND 1.24807f
C751 VDPWR.t23 VGND 0.003648f
C752 VDPWR.t56 VGND 0.003648f
C753 VDPWR.n66 VGND 0.007478f
C754 VDPWR.n67 VGND 0.061838f
C755 VDPWR.n68 VGND 0.019788f
C756 VDPWR.n69 VGND 0.044198f
C757 VDPWR.n70 VGND 0.049584f
C758 VDPWR.n71 VGND 0.049584f
C759 VDPWR.n72 VGND 0.3854f
C760 VDPWR.t32 VGND 0.152895f
C761 VDPWR.t42 VGND 0.106796f
C762 VDPWR.t26 VGND 0.059836f
C763 VDPWR.t28 VGND 0.072712f
C764 VDPWR.t36 VGND 0.119673f
C765 VDPWR.t24 VGND 0.119673f
C766 VDPWR.t30 VGND 0.154514f
C767 VDPWR.t59 VGND 0.039869f
C768 VDPWR.t58 VGND 0.039869f
C769 VDPWR.n73 VGND 0.054722f
C770 VDPWR.n74 VGND 0.010614f
C771 VDPWR.n75 VGND 0.039485f
C772 VDPWR.n76 VGND 0.046455f
C773 VDPWR.n77 VGND 0.044681f
C774 VDPWR.n78 VGND 0.022182f
C775 VDPWR.n79 VGND 0.049822f
C776 VDPWR.n80 VGND 0.209066f
C777 VDPWR.n81 VGND 0.100779f
C778 VDPWR.t40 VGND 0.217394f
C779 VDPWR.t22 VGND 0.173712f
C780 VDPWR.n82 VGND 0.150094f
C781 VDPWR.t55 VGND 0.299962f
C782 VDPWR.n83 VGND 0.326094f
C783 VDPWR.n84 VGND 0.049822f
C784 VDPWR.n85 VGND 0.045798f
C785 VDPWR.n86 VGND 0.024829f
C786 VDPWR.n87 VGND 0.029791f
C787 VDPWR.n88 VGND 0.019263f
C788 VDPWR.n89 VGND 0.649888f
C789 VDPWR.t50 VGND 0.001259f
C790 VDPWR.t43 VGND 0.001259f
C791 VDPWR.n90 VGND 0.002519f
C792 VDPWR.n91 VGND 0.003602f
C793 VDPWR.t33 VGND 0.001259f
C794 VDPWR.t46 VGND 0.001259f
C795 VDPWR.n92 VGND 0.002519f
C796 VDPWR.n93 VGND 0.003602f
C797 VDPWR.n94 VGND 0.076297f
C798 VDPWR.t29 VGND 0.001259f
C799 VDPWR.t45 VGND 0.001259f
C800 VDPWR.n95 VGND 0.002519f
C801 VDPWR.n96 VGND 0.003602f
C802 VDPWR.t47 VGND 0.001259f
C803 VDPWR.t37 VGND 0.001259f
C804 VDPWR.n97 VGND 0.002519f
C805 VDPWR.n98 VGND 0.003602f
C806 VDPWR.n99 VGND 0.117955f
C807 VDPWR.t48 VGND 0.001259f
C808 VDPWR.t31 VGND 0.001259f
C809 VDPWR.n100 VGND 0.002519f
C810 VDPWR.n101 VGND 0.003602f
C811 VDPWR.t25 VGND 0.001259f
C812 VDPWR.t49 VGND 0.001259f
C813 VDPWR.n102 VGND 0.002519f
C814 VDPWR.n103 VGND 0.003602f
C815 VDPWR.n104 VGND 0.024702f
C816 VDPWR.n105 VGND 0.074262f
C817 VDPWR.t27 VGND 0.003648f
C818 VDPWR.t41 VGND 0.003648f
C819 VDPWR.n106 VGND 0.007478f
C820 VDPWR.n107 VGND 0.020636f
C821 VDPWR.n108 VGND 0.03132f
C822 VDPWR.n109 VGND 0.456272f
C823 VDPWR.n110 VGND 0.633875f
C824 VDPWR.n111 VGND 0.014409f
C825 VDPWR.n112 VGND 0.061838f
C826 VDPWR.n113 VGND 0.019788f
C827 VDPWR.n114 VGND 0.044198f
C828 VDPWR.n115 VGND 0.049584f
C829 VDPWR.n116 VGND 0.049584f
C830 VDPWR.n117 VGND 0.3854f
C831 VDPWR.t9 VGND 0.152895f
C832 VDPWR.t5 VGND 0.106796f
C833 VDPWR.t7 VGND 0.059836f
C834 VDPWR.t13 VGND 0.072712f
C835 VDPWR.t0 VGND 0.119673f
C836 VDPWR.t15 VGND 0.119673f
C837 VDPWR.t3 VGND 0.154514f
C838 VDPWR.t61 VGND 0.039869f
C839 VDPWR.t60 VGND 0.039869f
C840 VDPWR.n118 VGND 0.054722f
C841 VDPWR.n119 VGND 0.010614f
C842 VDPWR.n120 VGND 0.039485f
C843 VDPWR.n121 VGND 0.046455f
C844 VDPWR.n122 VGND 0.044681f
C845 VDPWR.n123 VGND 0.022182f
C846 VDPWR.n124 VGND 0.049822f
C847 VDPWR.n125 VGND 0.209066f
C848 VDPWR.n126 VGND 0.100779f
C849 VDPWR.t53 VGND 0.217394f
C850 VDPWR.t38 VGND 0.173712f
C851 VDPWR.n127 VGND 0.150094f
C852 VDPWR.t34 VGND 0.299962f
C853 VDPWR.n128 VGND 0.326094f
C854 VDPWR.n129 VGND 0.049822f
C855 VDPWR.n130 VGND 0.045798f
C856 VDPWR.n131 VGND 0.024829f
C857 VDPWR.n132 VGND 0.029791f
C858 flash_0.x7.pos_en_b.n0 VGND 0.766491f
C859 flash_0.x7.pos_en_b.t6 VGND 0.932199f
C860 flash_0.x7.pos_en_b.t4 VGND 0.216253f
C861 flash_0.x7.pos_en_b.t5 VGND 0.216253f
C862 flash_0.x7.pos_en_b.t0 VGND 0.010089f
C863 flash_0.x7.pos_en_b.t1 VGND 0.010089f
C864 flash_0.x7.pos_en_b.t2 VGND 0.008975f
C865 flash_0.x7.pos_en_b.n1 VGND 0.032452f
C866 flash_0.x7.pos_en_b.t3 VGND 0.008975f
C867 flash_0.x4.dcgint.t0 VGND 0.016015f
C868 flash_0.x4.dcgint.t1 VGND 0.016015f
C869 flash_0.x4.dcgint.t2 VGND 0.016015f
C870 flash_0.x4.dcgint.t8 VGND 0.017561f
C871 flash_0.x4.dcgint.n0 VGND 0.05401f
C872 flash_0.x4.dcgint.t6 VGND 0.017266f
C873 flash_0.x4.dcgint.t9 VGND 0.355987f
C874 flash_0.x4.dcgint.t3 VGND 0.222316f
C875 flash_0.x4.dcgint.t5 VGND 0.280884f
C876 flash_0.x4.dcgint.t4 VGND 0.004616f
C877 flash_0.x4.dcgint.t10 VGND 0.004616f
C878 flash_0.x4.dcgint.n1 VGND 0.009325f
C879 flash_0.x4.dcgint.t7 VGND 0.004616f
C880 flash_0.x4.dcgint.t11 VGND 0.004616f
C881 flash_0.x4.dcgint.n2 VGND 0.009325f
C882 flash_0.x4.dcgint.n3 VGND 0.045712f
C883 flash_0.x4.dcgint.n4 VGND 0.233815f
C884 flash_0.x4.dcgint.n5 VGND 0.046322f
C885 flash_0.x4.dcgint.n6 VGND 0.34091f
C886 flash_0.x4.neg_mid_b.t10 VGND 0.828035f
C887 flash_0.x4.neg_mid_b.n0 VGND 0.140489f
C888 flash_0.x4.neg_mid_b.t1 VGND 0.007678f
C889 flash_0.x4.neg_mid_b.t2 VGND 0.007678f
C890 flash_0.x4.neg_mid_b.n1 VGND 0.015666f
C891 flash_0.x4.neg_mid_b.t0 VGND 0.02816f
C892 flash_0.x4.neg_mid_b.t7 VGND 0.067252f
C893 flash_0.x4.neg_mid_b.t8 VGND 0.122491f
C894 flash_0.x4.neg_mid_b.t12 VGND 0.067252f
C895 flash_0.x4.neg_mid_b.t14 VGND 0.122491f
C896 flash_0.x4.neg_mid_b.t11 VGND 0.067252f
C897 flash_0.x4.neg_mid_b.t13 VGND 0.122491f
C898 flash_0.x4.neg_mid_b.t3 VGND 0.007678f
C899 flash_0.x4.neg_mid_b.t6 VGND 0.007678f
C900 flash_0.x4.neg_mid_b.n2 VGND 0.015661f
C901 flash_0.x4.neg_mid_b.t4 VGND 0.02709f
C902 flash_0.x4.neg_mid_b.t9 VGND 0.085863f
C903 flash_0.x4.neg_mid_b.t5 VGND 0.027096f
C904 flash_0.x4.neg_en_b.n0 VGND 0.117521f
C905 flash_0.x4.neg_en_b.t0 VGND 0.036466f
C906 flash_0.x4.neg_en_b.t4 VGND 0.052338f
C907 flash_0.x4.neg_en_b.t8 VGND 0.051225f
C908 flash_0.x4.neg_en_b.t7 VGND 0.051225f
C909 flash_0.x4.neg_en_b.t5 VGND 0.051225f
C910 flash_0.x4.neg_en_b.t6 VGND 0.051201f
C911 flash_0.x4.neg_en_b.t9 VGND 0.051201f
C912 flash_0.x4.neg_en_b.t1 VGND 0.038945f
C913 flash_0.x4.neg_en_b.t2 VGND 0.032439f
C914 flash_0.x4.neg_en_b.t3 VGND 0.032439f
C915 ui_in[1].t17 VGND 0.038804f
C916 ui_in[1].n0 VGND 0.059281f
C917 ui_in[1].t10 VGND 0.038804f
C918 ui_in[1].n1 VGND 0.153087f
C919 ui_in[1].t12 VGND 0.038804f
C920 ui_in[1].n2 VGND 0.112696f
C921 ui_in[1].t13 VGND 0.038804f
C922 ui_in[1].n3 VGND 0.153087f
C923 ui_in[1].t15 VGND 0.038804f
C924 ui_in[1].n4 VGND 0.059281f
C925 ui_in[1].t2 VGND 0.038804f
C926 ui_in[1].n5 VGND 0.150815f
C927 ui_in[1].n6 VGND 0.419078f
C928 ui_in[1].t5 VGND 0.273311f
C929 ui_in[1].t0 VGND 0.285595f
C930 ui_in[1].n7 VGND 0.460636f
C931 ui_in[1].n8 VGND 0.339439f
C932 ui_in[1].t16 VGND 0.273311f
C933 ui_in[1].t14 VGND 0.285595f
C934 ui_in[1].n9 VGND 0.460636f
C935 ui_in[1].n10 VGND 0.233681f
C936 ui_in[1].n11 VGND 0.232247f
C937 ui_in[1].n12 VGND 0.130673f
C938 ui_in[1].n13 VGND 0.3368f
C939 ui_in[1].t7 VGND 0.228783f
C940 ui_in[1].t4 VGND 0.210357f
C941 ui_in[1].n14 VGND 0.322446f
C942 ui_in[1].n15 VGND 0.1233f
C943 ui_in[1].n16 VGND 0.166798f
C944 ui_in[1].t11 VGND 0.273311f
C945 ui_in[1].t8 VGND 0.285595f
C946 ui_in[1].n17 VGND 0.460636f
C947 ui_in[1].n18 VGND 0.229305f
C948 ui_in[1].n19 VGND 0.101954f
C949 ui_in[1].t9 VGND 0.273311f
C950 ui_in[1].t6 VGND 0.285595f
C951 ui_in[1].n20 VGND 0.460636f
C952 ui_in[1].n21 VGND 0.229305f
C953 ui_in[1].n22 VGND 0.102548f
C954 ui_in[1].n23 VGND 0.322167f
C955 ui_in[1].t3 VGND 0.228783f
C956 ui_in[1].t1 VGND 0.210357f
C957 ui_in[1].n24 VGND 0.322446f
C958 ui_in[1].n25 VGND 0.132755f
C959 ui_in[1].n26 VGND 0.521959f
C960 ui_in[1].n27 VGND 4.58386f
C961 ui_in[1].n28 VGND 0.52285f
C962 flash_0.x4.pos_mid_b.t1 VGND 0.019679f
C963 flash_0.x4.pos_mid_b.t2 VGND 0.019666f
C964 flash_0.x4.pos_mid_b.t8 VGND 0.055631f
C965 flash_0.x4.pos_mid_b.t7 VGND 0.055631f
C966 flash_0.x4.pos_mid_b.t4 VGND 0.055631f
C967 flash_0.x4.pos_mid_b.t3 VGND 0.055631f
C968 flash_0.x4.pos_mid_b.t6 VGND 0.055631f
C969 flash_0.x4.pos_mid_b.t5 VGND 0.055631f
C970 flash_0.x4.pos_mid_b.t0 VGND 0.020073f
C971 clk.t0 VGND 0.123904f
C972 clk.t1 VGND 0.116806f
C973 clk.n0 VGND 0.454326f
C974 clk.t2 VGND 0.123904f
C975 clk.t3 VGND 0.116806f
C976 clk.n1 VGND 0.454326f
C977 clk.n2 VGND 1.74152f
C978 clk.n3 VGND 4.1318f
C979 flash_0.x2.clkb.t1 VGND 0.011623f
C980 flash_0.x2.clkb.t0 VGND 0.018241f
C981 VAPWR.t6 VGND 0.003481f
C982 VAPWR.n0 VGND 0.025641f
C983 VAPWR.t1 VGND 0.003478f
C984 VAPWR.n1 VGND 0.034609f
C985 VAPWR.n2 VGND 0.04124f
C986 VAPWR.n3 VGND 0.025842f
C987 VAPWR.n4 VGND 0.045085f
C988 VAPWR.n5 VGND 0.148926f
C989 VAPWR.n6 VGND 0.050067f
C990 VAPWR.n7 VGND 0.050067f
C991 VAPWR.n8 VGND 0.022493f
C992 VAPWR.n9 VGND 0.022493f
C993 VAPWR.t8 VGND 0.010283f
C994 VAPWR.n10 VGND 0.022741f
C995 VAPWR.n11 VGND 0.130115f
C996 VAPWR.n12 VGND 0.130115f
C997 VAPWR.n13 VGND 0.183947f
C998 VAPWR.n14 VGND 0.049835f
C999 VAPWR.n15 VGND 0.022537f
C1000 VAPWR.n16 VGND 0.030498f
C1001 VAPWR.n17 VGND 0.022154f
C1002 VAPWR.n18 VGND 0.020469f
C1003 VAPWR.n19 VGND 0.030498f
C1004 VAPWR.n20 VGND 0.022537f
C1005 VAPWR.n21 VGND 0.048933f
C1006 VAPWR.n22 VGND 0.030426f
C1007 VAPWR.n23 VGND 0.022493f
C1008 VAPWR.n24 VGND 0.048933f
C1009 VAPWR.n25 VGND 0.190476f
C1010 VAPWR.n26 VGND 0.049075f
C1011 VAPWR.n27 VGND 0.183947f
C1012 VAPWR.n28 VGND 0.190476f
C1013 VAPWR.n29 VGND 0.183947f
C1014 VAPWR.n30 VGND 0.049075f
C1015 VAPWR.n31 VGND 0.016776f
C1016 VAPWR.n32 VGND 0.016833f
C1017 VAPWR.n33 VGND 0.022071f
C1018 VAPWR.n34 VGND 0.147307f
C1019 VAPWR.n35 VGND 0.020469f
C1020 VAPWR.n36 VGND 0.030498f
C1021 VAPWR.n37 VGND 0.022537f
C1022 VAPWR.n38 VGND 0.048933f
C1023 VAPWR.n39 VGND 0.030426f
C1024 VAPWR.n40 VGND 0.022493f
C1025 VAPWR.n41 VGND 0.049459f
C1026 VAPWR.n42 VGND 0.190476f
C1027 VAPWR.n43 VGND 0.049143f
C1028 VAPWR.n44 VGND 0.183947f
C1029 VAPWR.n45 VGND 0.190476f
C1030 VAPWR.n46 VGND 0.183947f
C1031 VAPWR.n47 VGND 0.049143f
C1032 VAPWR.n48 VGND 0.016776f
C1033 VAPWR.n49 VGND 0.016833f
C1034 VAPWR.n50 VGND 0.022071f
C1035 VAPWR.n51 VGND 0.034828f
C1036 VAPWR.n52 VGND 0.306925f
C1037 VAPWR.n53 VGND 0.083428f
C1038 VAPWR.n54 VGND 0.054859f
C1039 VAPWR.n55 VGND 0.073402f
C1040 VAPWR.n56 VGND 0.028091f
C1041 VAPWR.n57 VGND 0.022537f
C1042 VAPWR.n58 VGND 0.049832f
C1043 VAPWR.n59 VGND 0.15277f
C1044 VAPWR.n60 VGND 0.188825f
C1045 VAPWR.n61 VGND 0.135464f
C1046 VAPWR.n62 VGND 0.033985f
C1047 VAPWR.n63 VGND 0.015983f
C1048 VAPWR.t7 VGND 0.037542f
C1049 VAPWR.t5 VGND 0.343435f
C1050 VAPWR.t0 VGND 0.182547f
C1051 VAPWR.n64 VGND 0.142205f
C1052 VAPWR.n65 VGND 0.019665f
C1053 VAPWR.n66 VGND 0.026555f
C1054 VAPWR.n67 VGND 0.00647f
C1055 VAPWR.t13 VGND 0.010229f
C1056 VAPWR.n68 VGND 0.055175f
C1057 VAPWR.n69 VGND 0.059815f
C1058 VAPWR.n70 VGND 0.096071f
C1059 VAPWR.t16 VGND 0.003478f
C1060 VAPWR.n71 VGND 0.017733f
C1061 VAPWR.t10 VGND 0.003481f
C1062 VAPWR.n72 VGND 0.025711f
C1063 VAPWR.n73 VGND 0.045085f
C1064 VAPWR.n74 VGND 0.148926f
C1065 VAPWR.n75 VGND 0.050067f
C1066 VAPWR.n76 VGND 0.050067f
C1067 VAPWR.n77 VGND 0.022493f
C1068 VAPWR.n78 VGND 0.022493f
C1069 VAPWR.t12 VGND 0.010283f
C1070 VAPWR.n79 VGND 0.121994f
C1071 VAPWR.n80 VGND 0.01091f
C1072 VAPWR.n81 VGND 0.018798f
C1073 VAPWR.n82 VGND 0.011001f
C1074 VAPWR.n83 VGND 0.018798f
C1075 VAPWR.n84 VGND 0.085518f
C1076 VAPWR.t3 VGND 0.104521f
C1077 VAPWR.n87 VGND 0.085518f
C1078 VAPWR.t4 VGND 0.006509f
C1079 VAPWR.n88 VGND 0.040216f
C1080 VAPWR.n89 VGND 0.13191f
C1081 VAPWR.n90 VGND 0.065256f
C1082 VAPWR.n91 VGND 0.130115f
C1083 VAPWR.n92 VGND 0.130115f
C1084 VAPWR.n93 VGND 0.183947f
C1085 VAPWR.n94 VGND 0.049835f
C1086 VAPWR.n95 VGND 0.023894f
C1087 VAPWR.n96 VGND 0.094738f
C1088 VAPWR.t2 VGND 0.019586f
C1089 VAPWR.n97 VGND 0.006748f
C1090 VAPWR.n98 VGND 0.003219f
C1091 VAPWR.n99 VGND 0.057898f
C1092 VAPWR.n100 VGND 0.081102f
C1093 VAPWR.n101 VGND 0.023469f
C1094 VAPWR.n102 VGND 0.038288f
C1095 VAPWR.n103 VGND 0.030914f
C1096 VAPWR.n104 VGND 0.005625f
C1097 VAPWR.n105 VGND 0.027268f
C1098 VAPWR.n106 VGND 0.01091f
C1099 VAPWR.n107 VGND 0.011001f
C1100 VAPWR.n108 VGND 0.018067f
C1101 VAPWR.n109 VGND 0.022537f
C1102 VAPWR.n110 VGND 0.049832f
C1103 VAPWR.n111 VGND 0.15277f
C1104 VAPWR.n112 VGND 0.188825f
C1105 VAPWR.n113 VGND 0.135464f
C1106 VAPWR.n114 VGND 0.033985f
C1107 VAPWR.n115 VGND 0.015983f
C1108 VAPWR.t11 VGND 0.037542f
C1109 VAPWR.t9 VGND 0.343435f
C1110 VAPWR.t15 VGND 0.182547f
C1111 VAPWR.n116 VGND 0.142205f
C1112 VAPWR.n117 VGND 0.019665f
C1113 VAPWR.n118 VGND 0.026555f
C1114 VAPWR.n119 VGND 0.018775f
C1115 VAPWR.t14 VGND 0.010259f
C1116 VAPWR.n120 VGND 0.094854f
C1117 VAPWR.n121 VGND 0.11419f
C1118 VAPWR.n122 VGND 0.018245f
C1119 VAPWR.n123 VGND 1.0575f
C1120 VAPWR.n124 VGND 0.521869f
C1121 VAPWR.n125 VGND 7.2806f
C1122 VAPWR.n126 VGND 40.983803f
C1123 flash_0.x7.VPRGPOS.t27 VGND 0.001388f
C1124 flash_0.x7.VPRGPOS.t16 VGND 0.040919f
C1125 flash_0.x7.VPRGPOS.t11 VGND 0.025964f
C1126 flash_0.x7.VPRGPOS.t12 VGND 0.025964f
C1127 flash_0.x7.VPRGPOS.t15 VGND 0.025964f
C1128 flash_0.x7.VPRGPOS.t13 VGND 0.025471f
C1129 flash_0.x7.VPRGPOS.t23 VGND 0.111581f
C1130 flash_0.x7.VPRGPOS.t14 VGND 0.043055f
C1131 flash_0.x7.VPRGPOS.n0 VGND 0.00573f
C1132 flash_0.x7.VPRGPOS.t24 VGND 0.001388f
C1133 flash_0.x7.VPRGPOS.t30 VGND 0.001388f
C1134 flash_0.x7.VPRGPOS.t10 VGND 0.002773f
C1135 flash_0.x7.VPRGPOS.t1 VGND 0.001483f
C1136 flash_0.x7.VPRGPOS.n1 VGND 0.021758f
C1137 flash_0.x7.VPRGPOS.n2 VGND 0.021822f
C1138 flash_0.x7.VPRGPOS.n4 VGND 0.037489f
C1139 flash_0.x7.VPRGPOS.n5 VGND 0.022319f
C1140 flash_0.x7.VPRGPOS.n6 VGND 0.256188f
C1141 flash_0.x7.VPRGPOS.t0 VGND 0.411174f
C1142 flash_0.x7.VPRGPOS.n8 VGND 0.037489f
C1143 flash_0.x7.VPRGPOS.n9 VGND 0.256188f
C1144 flash_0.x7.VPRGPOS.n10 VGND 0.012323f
C1145 flash_0.x7.VPRGPOS.n11 VGND 0.01234f
C1146 flash_0.x7.VPRGPOS.n12 VGND 0.026121f
C1147 flash_0.x7.VPRGPOS.t18 VGND 0.001388f
C1148 flash_0.x7.VPRGPOS.t7 VGND 3.92e-19
C1149 flash_0.x7.VPRGPOS.t5 VGND 3.92e-19
C1150 flash_0.x7.VPRGPOS.n13 VGND 8.05e-19
C1151 flash_0.x7.VPRGPOS.t32 VGND 3.92e-19
C1152 flash_0.x7.VPRGPOS.t9 VGND 3.92e-19
C1153 flash_0.x7.VPRGPOS.n14 VGND 8.05e-19
C1154 flash_0.x7.VPRGPOS.t20 VGND 0.001388f
C1155 flash_0.x7.VPRGPOS.t17 VGND 0.040919f
C1156 flash_0.x7.VPRGPOS.t6 VGND 0.025964f
C1157 flash_0.x7.VPRGPOS.t4 VGND 0.025964f
C1158 flash_0.x7.VPRGPOS.t21 VGND 0.025964f
C1159 flash_0.x7.VPRGPOS.t8 VGND 0.025471f
C1160 flash_0.x7.VPRGPOS.t2 VGND 0.111581f
C1161 flash_0.x7.VPRGPOS.t19 VGND 0.043055f
C1162 flash_0.x7.VPRGPOS.n15 VGND 0.00573f
C1163 flash_0.x7.VPRGPOS.t31 VGND 0.001388f
C1164 flash_0.x7.VPRGPOS.t3 VGND 0.001388f
C1165 flash_0.x7.VPRGPOS.n16 VGND 0.098365f
C1166 flash_0.x7.VPRGPOS.n17 VGND 1.69352f
C1167 flash_0.x7.VPRGPOS.t25 VGND 0.001388f
C1168 flash_0.x7.VPRGPOS.t26 VGND 3.92e-19
C1169 flash_0.x7.VPRGPOS.t22 VGND 3.92e-19
C1170 flash_0.x7.VPRGPOS.n18 VGND 8.05e-19
C1171 flash_0.x7.VPRGPOS.t28 VGND 3.92e-19
C1172 flash_0.x7.VPRGPOS.t29 VGND 3.92e-19
C1173 flash_0.x7.VPRGPOS.n19 VGND 8.05e-19
C1174 flash_0.x7.pos_mid_b.t2 VGND 0.020534f
C1175 flash_0.x7.pos_mid_b.t0 VGND 0.020521f
C1176 flash_0.x7.pos_mid_b.t4 VGND 0.020534f
C1177 flash_0.x7.pos_mid_b.t1 VGND 0.020521f
C1178 flash_0.x7.pos_mid_b.t3 VGND 0.020946f
C1179 flash_0.x7.pos_mid_b.t9 VGND 0.05805f
C1180 flash_0.x7.pos_mid_b.t10 VGND 0.05805f
C1181 flash_0.x7.pos_mid_b.t8 VGND 0.05805f
C1182 flash_0.x7.pos_mid_b.t5 VGND 0.05805f
C1183 flash_0.x7.pos_mid_b.t6 VGND 0.05805f
C1184 flash_0.x7.pos_mid_b.t7 VGND 0.05805f
.ends

