* NGSPICE file created from vprog_controller.ext - technology: sky130A
.subckt vprog_controller pos_en neg_en VOUT VDPWR VGND VPRGPOS VPRGNEG
X0 pos_mid_b.t2 pos_en.t0 VGND.t8 VGND.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X1 VOUT.t3 neg_mid_b dcgint dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X2 VDPWR pos_en.t1 pos_en_b.t2 VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X3 VOUT.t7 VDPWR vintp VPRGPOS.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X4 dcgint neg_mid_b VOUT.t2 dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X5 pos_mid_b pos_en.t0 VGND.t7 VGND.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X6 vintp pos_mid_b.t4 VPRGPOS.t10 VPRGPOS.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X7 neg_en_b.t1 neg_en.t0 VGND.t21 VGND.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X8 VPRGPOS pos_mid_b vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X9 VOUT.t1 neg_mid_b dcgint dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X10 dcgint neg_mid_b VOUT.t0 dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X11 neg_mid neg_en.t1 VDPWR.t12 VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X12 pos_mid pos_en_b.t3 VGND.t19 VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X13 neg_en_b neg_en.t2 VDPWR.t15 VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=3
X14 VDPWR neg_en_b neg_mid_b VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X15 VDPWR.t13 neg_en_b.t3 neg_mid_b VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X16 vintp pos_mid_b.t5 VPRGPOS.t8 VPRGPOS.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X17 a_2408_n3852# neg_mid_b VPRGNEG.t5 VPRGNEG.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X18 VDPWR.t10 neg_en_b.t4 neg_mid_b VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X19 vintp VDPWR VOUT.t6 VPRGPOS.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X20 pos_mid pos_en_b.t3 VGND.t18 VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X21 neg_mid neg_en.t3 VDPWR.t0 VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X22 neg_mid neg_en.t4 VDPWR.t8 VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X23 VOUT VDPWR vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X24 VGND.t11 pos_en_b.t4 pos_mid VGND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X25 pos_en_b.t1 pos_en.t2 VGND.t5 VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X26 a_2408_n3852# neg_mid_b VPRGNEG.t3 VPRGNEG.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=3
X27 vintp VDPWR VOUT.t5 VPRGPOS.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X28 VGND.t10 pos_en_b.t4 pos_mid VGND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X29 pos_en_b pos_en.t3 VDPWR VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.21 ps=1.34 w=0.5 l=3
X30 VPRGPOS pos_mid_b vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X31 VGND.t20 neg_en.t5 neg_en_b.t0 VGND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X32 vintp pos_mid_b.t6 VPRGPOS.t6 VPRGPOS.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X33 dcgint pos_en_b.t5 VGND.t17 VGND.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X34 VDPWR neg_en neg_mid VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.135 ps=1.54 w=0.5 l=0.5
X35 VDPWR.t6 neg_en.t6 neg_en_b.t2 VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X36 VDPWR.t14 neg_en.t7 neg_mid VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X37 dcgint pos_en_b.t5 VGND.t15 VGND.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X38 VPRGPOS.t1 pos_mid pos_mid_b.t3 VPRGPOS.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X39 neg_mid_b neg_mid VPRGNEG.t6 VPRGNEG.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.21 ps=1.34 w=0.5 l=1
X40 neg_mid_b neg_en_b.t5 VDPWR.t7 VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X41 neg_mid_b neg_en_b.t6 VDPWR.t9 VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X42 VPRGNEG.t1 neg_mid_b neg_mid VPRGNEG.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.145 ps=1.58 w=0.5 l=1
X43 VOUT VDPWR vintp VPRGPOS sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.5
X44 vintp VDPWR VOUT.t4 VPRGPOS.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X45 dcgint neg_mid_b VOUT dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X46 VGND.t3 pos_en.t4 pos_mid_b.t1 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X47 dcgint pos_en_b.t5 VGND.t13 VGND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X48 VOUT VDPWR a_2408_n3852# VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X49 VPRGPOS.t4 pos_mid_b.t7 pos_mid VPRGPOS.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.135 ps=1.54 w=0.5 l=3
X50 VGND.t2 pos_en.t4 pos_mid_b.t0 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X51 VOUT VDPWR a_2408_n3852# VPRGNEG sky130_fd_pr__nfet_g5v0d10v5 ad=0.135 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=3
X52 VPRGPOS.t3 pos_mid_b.t8 vintp VPRGPOS.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X53 neg_mid_b neg_en_b.t7 VDPWR.t5 VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X54 dcgint neg_mid_b VOUT dcgint sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X55 VGND.t1 pos_en.t5 pos_en_b.t0 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.34 as=0.135 ps=1.54 w=0.5 l=3
X56 VDPWR.t11 neg_en.t8 neg_mid VDPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
C0 VDPWR VPRGNEG 6.45435f
C1 neg_mid_b dcgint 2.14914f
C2 neg_en VDPWR 2.05821f
C3 neg_en neg_en_b 3.01537f
C4 VPRGNEG neg_mid_b 2.17163f
C5 pos_mid_b VPRGPOS 2.22569f
C6 pos_en_b pos_en 2.34221f
R0 pos_en.n0 pos_en 123.99
R1 pos_en.t4 pos_en.n3 114.805
R2 pos_en pos_en.n0 50.8126
R3 pos_en.n0 pos_en 29.418
R4 pos_en.n0 pos_en 29.418
R5 pos_en.n0 pos_en.t4 24.0464
R6 pos_en.n0 pos_en.n2 19.0005
R7 pos_en.n0 pos_en.n1 19.0005
R8 pos_en pos_en.t0 19.0005
R9 pos_en.n2 pos_en.t5 12.0505
R10 pos_en.n2 pos_en.t1 12.0505
R11 pos_en.n1 pos_en.t2 12.0505
R12 pos_en.n1 pos_en.t3 12.0505
R13 VGND.n8 VGND.n1 3014.19
R14 VGND.t16 VGND.n9 16658.8
R15 VGND.t9 VGND.t4 4288.33
R16 VGND.t4 VGND.t0 4288.33
R17 VGND.t6 VGND.n8 3495.43
R18 VGND.n9 VGND.n1 3250.9
R19 VGND.n9 VGND.t6 2825.38
R20 VGND.t0 VGND 2659.27
R21 VGND.n8 VGND.t9 792.894
R22 VGND.t14 VGND.t16 712.963
R23 VGND.n10 VGND.t12 444.753
R24 VGND.n10 VGND.t14 268.211
R25 VGND VGND.t17 230.898
R26 VGND VGND.t15 230.898
R27 VGND.n0 VGND.t13 218.06
R28 VGND.n1 VGND 1.75967
R29 VGND VGND.n7 97.1505
R30 VGND VGND.n4 97.1505
R31 VGND VGND.n5 97.1505
R32 VGND VGND.n2 97.1505
R33 VGND VGND.n6 97.1505
R34 VGND VGND.n3 97.1505
R35 VGND.n7 VGND.t19 95.7605
R36 VGND.n7 VGND.t3 95.7605
R37 VGND.n4 VGND.t8 95.7605
R38 VGND.n4 VGND.t11 95.7605
R39 VGND.n5 VGND.t18 95.7605
R40 VGND.n5 VGND.t2 95.7605
R41 VGND.n2 VGND.t7 95.7605
R42 VGND.n2 VGND.t10 95.7605
R43 VGND.n6 VGND.t5 95.7605
R44 VGND.n6 VGND.t1 95.7605
R45 VGND.n3 VGND.t21 95.7605
R46 VGND.n3 VGND.t20 95.7605
R47 VGND.n10 VGND 73.8569
R48 VGND VGND.n0 23.4721
R49 pos_mid_b pos_mid_b.t3 649.691
R50 pos_mid_b pos_mid_b.t1 227.361
R51 pos_mid_b pos_mid_b.t0 227.361
R52 pos_mid_b pos_mid_b.t2 227.361
R53 pos_mid_b pos_mid_b.t4 216.731
R54 pos_mid_b pos_mid_b.n0 216.731
R55 pos_mid_b pos_mid_b.t6 216.731
R56 pos_mid_b pos_mid_b.t8 216.731
R57 pos_mid_b pos_mid_b.t5 216.731
R58 pos_mid_b pos_mid_b.n1 216.731
R59 pos_mid_b pos_mid_b.t7 38.3118
R60 VOUT VOUT.t6 649.691
R61 VOUT VOUT.t4 649.691
R62 VOUT VOUT.n2 594.383
R63 VOUT VOUT.n1 594.301
R64 VOUT VOUT.n3 594.301
R65 VOUT.n1 VOUT.t5 55.3905
R66 VOUT.n1 VOUT.t7 55.3905
R67 VOUT.n3 VOUT.t2 55.3905
R68 VOUT.n3 VOUT.t3 55.3905
R69 VOUT.n2 VOUT.t0 55.3905
R70 VOUT.n2 VOUT.t1 55.3905
R71 VOUT VOUT.n0 16.7521
R72 pos_en_b pos_en_b.t2 640.39
R73 pos_en_b.n0 pos_en_b.t0 247.151
R74 pos_en_b.n1 pos_en_b.t1 247.151
R75 pos_en_b.n0 pos_en_b.t5 65.4032
R76 pos_en_b.t5 pos_en_b 56.2429
R77 pos_en_b.t5 pos_en_b 56.2429
R78 pos_en_b.n0 pos_en_b 50.8126
R79 pos_en_b.n0 pos_en_b 50.8126
R80 pos_en_b pos_en_b.n1 29.0914
R81 pos_en_b.n0 pos_en_b 29.0914
R82 pos_en_b.n1 pos_en_b.n0 28.2591
R83 pos_en_b.n0 pos_en_b.t3 27.4355
R84 pos_en_b.n0 pos_en_b.t4 27.4355
R85 VDPWR.n9 VDPWR.t0 640.39
R86 VDPWR.n8 VDPWR.n7 585
R87 VDPWR.n4 VDPWR.n3 585
R88 VDPWR.n6 VDPWR.n5 585
R89 VDPWR.n2 VDPWR.n1 585
R90 VDPWR.n12 VDPWR.n11 585
R91 VDPWR VDPWR.n0 297.151
R92 VDPWR.n0 VDPWR.t15 160.44
R93 VDPWR.n0 VDPWR.t6 160.44
R94 VDPWR.n7 VDPWR.t12 55.3905
R95 VDPWR.n7 VDPWR.t10 55.3905
R96 VDPWR.n3 VDPWR.t9 55.3905
R97 VDPWR.n3 VDPWR.t14 55.3905
R98 VDPWR.n5 VDPWR.t5 55.3905
R99 VDPWR.n5 VDPWR.t11 55.3905
R100 VDPWR.n1 VDPWR.t8 55.3905
R101 VDPWR.n1 VDPWR.t13 55.3905
R102 VDPWR.n11 VDPWR.t7 55.3905
R103 VDPWR.n11 VDPWR.n10 32.4705
R104 VDPWR VDPWR.n4 16.4381
R105 VDPWR.n8 VDPWR 14.3064
R106 VDPWR.n4 VDPWR 14.3064
R107 VDPWR.n9 VDPWR 14.3064
R108 VDPWR.n6 VDPWR 14.3064
R109 VDPWR.n2 VDPWR 14.3064
R110 VDPWR VDPWR.n12 14.3064
R111 VDPWR.n12 VDPWR 13.8019
R112 VDPWR VDPWR.n8 13.8019
R113 VDPWR VDPWR.n9 13.8019
R114 VDPWR VDPWR.n6 13.8019
R115 VDPWR VDPWR.n2 13.8019
R116 VPRGPOS.t9 VPRGPOS.t0 809.375
R117 VPRGPOS VPRGPOS.t4 649.691
R118 VPRGPOS VPRGPOS.t1 649.691
R119 VPRGPOS VPRGPOS.t10 649.691
R120 VPRGPOS VPRGPOS.t6 649.691
R121 VPRGPOS VPRGPOS.n1 594.301
R122 VPRGPOS.t9 VPRGPOS.t5 484.375
R123 VPRGPOS.t2 VPRGPOS.t7 246.875
R124 VPRGPOS.t5 VPRGPOS.t2 246.875
R125 VPRGPOS.n1 VPRGPOS.t8 55.3905
R126 VPRGPOS.n1 VPRGPOS.t3 55.3905
R127 VPRGPOS VPRGPOS.n0 43.6711
R128 VPRGPOS VPRGPOS.t9 27.4882
R129 neg_en neg_en.n2 207.43
R130 neg_en neg_en.t1 207.43
R131 neg_en neg_en.t7 207.43
R132 neg_en neg_en.t3 207.43
R133 neg_en neg_en.t8 207.43
R134 neg_en neg_en.t4 207.43
R135 neg_en neg_en.n0 25.4765
R136 neg_en neg_en.n1 19.0005
R137 neg_en.n0 neg_en.t5 12.0505
R138 neg_en.n0 neg_en.t6 12.0505
R139 neg_en.n1 neg_en.t0 12.0505
R140 neg_en.n1 neg_en.t2 12.0505
R141 neg_en_b neg_en_b.t2 640.39
R142 neg_en_b neg_en_b.t0 247.151
R143 neg_en_b.n1 neg_en_b.t1 247.151
R144 neg_en_b neg_en_b.t6 211.017
R145 neg_en_b neg_en_b.t5 208.394
R146 neg_en_b neg_en_b.t4 208.394
R147 neg_en_b neg_en_b.n0 207.43
R148 neg_en_b neg_en_b.t7 207.43
R149 neg_en_b neg_en_b.t3 207.43
R150 neg_en_b.n1 neg_en_b 50.3013
R151 neg_en_b neg_en_b.n1 29.0914
R152 VPRGNEG.n9 VPRGNEG.n6 6482.77
R153 VPRGNEG.n9 VPRGNEG.n2 6482.77
R154 VPRGNEG.n7 VPRGNEG.n2 6482.77
R155 VPRGNEG.n7 VPRGNEG.n6 6482.77
R156 VPRGNEG.t0 VPRGNEG.n8 565.485
R157 VPRGNEG.t4 VPRGNEG.t2 565.485
R158 VPRGNEG.n9 VPRGNEG.t0 530.141
R159 VPRGNEG.t2 VPRGNEG.n7 406.274
R160 VPRGNEG.n5 VPRGNEG.n4 287.248
R161 VPRGNEG.n5 VPRGNEG.n1 263.668
R162 VPRGNEG VPRGNEG.t5 227.361
R163 VPRGNEG.n0 VPRGNEG.t3 218.06
R164 VPRGNEG VPRGNEG.n10 164.915
R165 VPRGNEG.n8 VPRGNEG.t4 123.868
R166 VPRGNEG.n3 VPRGNEG.t6 95.7605
R167 VPRGNEG.n3 VPRGNEG.t1 95.7605
R168 VPRGNEG.n10 VPRGNEG.n4 95.2476
R169 VPRGNEG VPRGNEG.n3 92.5005
R170 VPRGNEG VPRGNEG.n1 87.7182
R171 VPRGNEG.n6 VPRGNEG.n5 58.5005
R172 VPRGNEG.n8 VPRGNEG.n6 58.5005
R173 VPRGNEG VPRGNEG.n2 58.5005
R174 VPRGNEG.n8 VPRGNEG.n2 58.5005
R175 VPRGNEG.n10 VPRGNEG.n9 26.5914
R176 VPRGNEG.n7 VPRGNEG.n1 26.5914
R177 VPRGNEG.n4 VPRGNEG 17.3454
R178 VPRGNEG.n0 VPRGNEG.n11 14.3064
R179 VPRGNEG VPRGNEG.n0 12.4535
C7 VDPWR VGND 24.64152f
C8 neg_en VGND 6.27242f
C9 pos_en VGND 7.18439f
C10 VPRGPOS VGND 4.48067f
C11 neg_en_b VGND 3.149f $ **FLOATING
C12 pos_en_b VGND 7.73169f $ **FLOATING
C13 neg_mid_b VGND 2.03401f $ **FLOATING
C14 pos_mid_b VGND 3.4665f $ **FLOATING
C15 dcgint VGND 2.90806f $ **FLOATING
.ends
