magic
tech sky130A
magscale 1 2
timestamp 1739996772
<< error_p >>
rect -519 267 519 553
rect -519 -267 -233 267
rect -29 117 29 123
rect -29 83 -17 117
rect -29 77 29 83
rect -29 -83 29 -77
rect -29 -117 -17 -83
rect -29 -123 29 -117
rect 233 -267 519 267
rect -519 -553 519 -267
<< dnwell >>
rect -439 -473 439 473
<< pwell >>
rect -221 -255 221 255
<< nsonos >>
rect -22 -45 22 45
<< ndiff >>
rect -83 33 -22 45
rect -83 -33 -71 33
rect -37 -33 -22 33
rect -83 -45 -22 -33
rect 22 33 83 45
rect 22 -33 37 33
rect 71 -33 83 33
rect 22 -45 83 -33
<< ndiffc >>
rect -71 -33 -37 33
rect 37 -33 71 33
<< psubdiff >>
rect -185 185 -89 219
rect 89 185 185 219
rect -185 123 -151 185
rect 151 123 185 185
rect -185 -185 -151 -123
rect 151 -185 185 -123
rect -185 -219 -89 -185
rect 89 -219 185 -185
<< psubdiffcont >>
rect -89 185 89 219
rect -185 -123 -151 123
rect 151 -123 185 123
rect -89 -219 89 -185
<< poly >>
rect -33 117 33 133
rect -33 83 -17 117
rect 17 83 33 117
rect -33 67 33 83
rect -22 45 22 67
rect -22 -67 22 -45
rect -33 -83 33 -67
rect -33 -117 -17 -83
rect 17 -117 33 -83
rect -33 -133 33 -117
<< polycont >>
rect -17 83 17 117
rect -17 -117 17 -83
<< locali >>
rect -185 185 -89 219
rect 89 185 185 219
rect -185 123 -151 185
rect 151 123 185 185
rect -33 83 -17 117
rect 17 83 33 117
rect -71 33 -37 49
rect -71 -49 -37 -33
rect 37 33 71 49
rect 37 -49 71 -33
rect -33 -117 -17 -83
rect 17 -117 33 -83
rect -185 -185 -151 -123
rect 151 -185 185 -123
rect -185 -219 -89 -185
rect 89 -219 185 -185
<< viali >>
rect -17 83 17 117
rect -71 -33 -37 33
rect 37 -33 71 33
rect -17 -117 17 -83
<< metal1 >>
rect -29 117 29 123
rect -29 83 -17 117
rect 17 83 29 117
rect -29 77 29 83
rect -77 33 -31 45
rect -77 -33 -71 33
rect -37 -33 -31 33
rect -77 -45 -31 -33
rect 31 33 77 45
rect 31 -33 37 33
rect 71 -33 77 33
rect 31 -45 77 -33
rect -29 -83 29 -77
rect -29 -117 -17 -83
rect 17 -117 29 -83
rect -29 -123 29 -117
<< properties >>
string FIXED_BBOX -168 -202 168 202
string gencell sky130_fd_bs_flash__special_sonosfet_star
string library sky130
string parameters w 0.45 l 0.22 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
